module ttsimon (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire net4;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire net3;
 wire net2;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire net108;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire net107;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire net106;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire net105;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire net104;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire net103;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire net102;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire net101;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire net100;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire net99;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire net98;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire net97;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire net96;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire _0662_;
 wire _0663_;
 wire net91;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire _0669_;
 wire _0670_;
 wire net85;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire net84;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire net83;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire net82;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire net81;
 wire _0708_;
 wire net80;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire net79;
 wire _0738_;
 wire _0739_;
 wire net78;
 wire net77;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire net76;
 wire net75;
 wire _0748_;
 wire _0749_;
 wire net74;
 wire net73;
 wire net72;
 wire _0753_;
 wire _0754_;
 wire net71;
 wire net70;
 wire net69;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire net68;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire net67;
 wire _0784_;
 wire _0785_;
 wire net66;
 wire _0787_;
 wire _0788_;
 wire net65;
 wire net64;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire net63;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire net62;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire net61;
 wire _0814_;
 wire net60;
 wire _0816_;
 wire net59;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire net58;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire net57;
 wire net56;
 wire net55;
 wire _0830_;
 wire net54;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire net53;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire net52;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire net51;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire net50;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire net49;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire net48;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire net47;
 wire net46;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire net45;
 wire _0900_;
 wire _0901_;
 wire net44;
 wire net43;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire net42;
 wire net41;
 wire _0913_;
 wire net40;
 wire _0915_;
 wire net39;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire net38;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire net37;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire net36;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire net35;
 wire _0963_;
 wire _0964_;
 wire net34;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire net33;
 wire net32;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire net31;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire net30;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire net29;
 wire _1029_;
 wire _1030_;
 wire net28;
 wire _1032_;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire net23;
 wire _1041_;
 wire net22;
 wire _1043_;
 wire net21;
 wire net20;
 wire _1046_;
 wire net19;
 wire net18;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire net17;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire net16;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire net15;
 wire net14;
 wire _1067_;
 wire net13;
 wire _1069_;
 wire net12;
 wire _1071_;
 wire net11;
 wire net10;
 wire _1074_;
 wire _1075_;
 wire net9;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire net8;
 wire _1086_;
 wire _1087_;
 wire net7;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire net6;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire net5;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire net1;
 wire \simon1.millis_counter[0] ;
 wire \simon1.millis_counter[1] ;
 wire \simon1.millis_counter[2] ;
 wire \simon1.millis_counter[3] ;
 wire \simon1.millis_counter[4] ;
 wire \simon1.millis_counter[5] ;
 wire \simon1.millis_counter[6] ;
 wire \simon1.millis_counter[7] ;
 wire \simon1.millis_counter[8] ;
 wire \simon1.millis_counter[9] ;
 wire \simon1.next_random[0] ;
 wire \simon1.next_random[1] ;
 wire \simon1.play1.freq[0] ;
 wire \simon1.play1.freq[1] ;
 wire \simon1.play1.freq[2] ;
 wire \simon1.play1.freq[3] ;
 wire \simon1.play1.freq[4] ;
 wire \simon1.play1.freq[5] ;
 wire \simon1.play1.freq[6] ;
 wire \simon1.play1.freq[7] ;
 wire \simon1.play1.freq[8] ;
 wire \simon1.play1.freq[9] ;
 wire \simon1.play1.tick_counter[0] ;
 wire \simon1.play1.tick_counter[10] ;
 wire \simon1.play1.tick_counter[11] ;
 wire \simon1.play1.tick_counter[12] ;
 wire \simon1.play1.tick_counter[13] ;
 wire \simon1.play1.tick_counter[14] ;
 wire \simon1.play1.tick_counter[15] ;
 wire \simon1.play1.tick_counter[16] ;
 wire \simon1.play1.tick_counter[17] ;
 wire \simon1.play1.tick_counter[18] ;
 wire \simon1.play1.tick_counter[19] ;
 wire \simon1.play1.tick_counter[1] ;
 wire \simon1.play1.tick_counter[20] ;
 wire \simon1.play1.tick_counter[21] ;
 wire \simon1.play1.tick_counter[22] ;
 wire \simon1.play1.tick_counter[23] ;
 wire \simon1.play1.tick_counter[24] ;
 wire \simon1.play1.tick_counter[25] ;
 wire \simon1.play1.tick_counter[26] ;
 wire \simon1.play1.tick_counter[27] ;
 wire \simon1.play1.tick_counter[28] ;
 wire \simon1.play1.tick_counter[29] ;
 wire \simon1.play1.tick_counter[2] ;
 wire \simon1.play1.tick_counter[30] ;
 wire \simon1.play1.tick_counter[31] ;
 wire \simon1.play1.tick_counter[3] ;
 wire \simon1.play1.tick_counter[4] ;
 wire \simon1.play1.tick_counter[5] ;
 wire \simon1.play1.tick_counter[6] ;
 wire \simon1.play1.tick_counter[7] ;
 wire \simon1.play1.tick_counter[8] ;
 wire \simon1.play1.tick_counter[9] ;
 wire \simon1.score1.active_digit ;
 wire \simon1.score1.ena ;
 wire \simon1.score1.inc ;
 wire \simon1.score1.ones[0] ;
 wire \simon1.score1.ones[1] ;
 wire \simon1.score1.ones[2] ;
 wire \simon1.score1.ones[3] ;
 wire \simon1.score1.tens[0] ;
 wire \simon1.score1.tens[1] ;
 wire \simon1.score1.tens[2] ;
 wire \simon1.score1.tens[3] ;
 wire \simon1.score_rst ;
 wire \simon1.seq[0][0] ;
 wire \simon1.seq[0][1] ;
 wire \simon1.seq[10][0] ;
 wire \simon1.seq[10][1] ;
 wire \simon1.seq[11][0] ;
 wire \simon1.seq[11][1] ;
 wire \simon1.seq[12][0] ;
 wire \simon1.seq[12][1] ;
 wire \simon1.seq[13][0] ;
 wire \simon1.seq[13][1] ;
 wire \simon1.seq[14][0] ;
 wire \simon1.seq[14][1] ;
 wire \simon1.seq[15][0] ;
 wire \simon1.seq[15][1] ;
 wire \simon1.seq[16][0] ;
 wire \simon1.seq[16][1] ;
 wire \simon1.seq[17][0] ;
 wire \simon1.seq[17][1] ;
 wire \simon1.seq[18][0] ;
 wire \simon1.seq[18][1] ;
 wire \simon1.seq[19][0] ;
 wire \simon1.seq[19][1] ;
 wire \simon1.seq[1][0] ;
 wire \simon1.seq[1][1] ;
 wire \simon1.seq[20][0] ;
 wire \simon1.seq[20][1] ;
 wire \simon1.seq[21][0] ;
 wire \simon1.seq[21][1] ;
 wire \simon1.seq[22][0] ;
 wire \simon1.seq[22][1] ;
 wire \simon1.seq[23][0] ;
 wire \simon1.seq[23][1] ;
 wire \simon1.seq[24][0] ;
 wire \simon1.seq[24][1] ;
 wire \simon1.seq[25][0] ;
 wire \simon1.seq[25][1] ;
 wire \simon1.seq[26][0] ;
 wire \simon1.seq[26][1] ;
 wire \simon1.seq[27][0] ;
 wire \simon1.seq[27][1] ;
 wire \simon1.seq[28][0] ;
 wire \simon1.seq[28][1] ;
 wire \simon1.seq[29][0] ;
 wire \simon1.seq[29][1] ;
 wire \simon1.seq[2][0] ;
 wire \simon1.seq[2][1] ;
 wire \simon1.seq[30][0] ;
 wire \simon1.seq[30][1] ;
 wire \simon1.seq[31][0] ;
 wire \simon1.seq[31][1] ;
 wire \simon1.seq[3][0] ;
 wire \simon1.seq[3][1] ;
 wire \simon1.seq[4][0] ;
 wire \simon1.seq[4][1] ;
 wire \simon1.seq[5][0] ;
 wire \simon1.seq[5][1] ;
 wire \simon1.seq[6][0] ;
 wire \simon1.seq[6][1] ;
 wire \simon1.seq[7][0] ;
 wire \simon1.seq[7][1] ;
 wire \simon1.seq[8][0] ;
 wire \simon1.seq[8][1] ;
 wire \simon1.seq[9][0] ;
 wire \simon1.seq[9][1] ;
 wire \simon1.seq_counter[0] ;
 wire \simon1.seq_counter[1] ;
 wire \simon1.seq_counter[2] ;
 wire \simon1.seq_counter[3] ;
 wire \simon1.seq_counter[4] ;
 wire \simon1.seq_length[0] ;
 wire \simon1.seq_length[1] ;
 wire \simon1.seq_length[2] ;
 wire \simon1.seq_length[3] ;
 wire \simon1.seq_length[4] ;
 wire \simon1.state[0] ;
 wire \simon1.state[1] ;
 wire \simon1.state[2] ;
 wire \simon1.state[3] ;
 wire \simon1.state[4] ;
 wire \simon1.state[5] ;
 wire \simon1.state[6] ;
 wire \simon1.state[7] ;
 wire \simon1.tick_counter[0] ;
 wire \simon1.tick_counter[10] ;
 wire \simon1.tick_counter[11] ;
 wire \simon1.tick_counter[12] ;
 wire \simon1.tick_counter[13] ;
 wire \simon1.tick_counter[14] ;
 wire \simon1.tick_counter[15] ;
 wire \simon1.tick_counter[1] ;
 wire \simon1.tick_counter[2] ;
 wire \simon1.tick_counter[3] ;
 wire \simon1.tick_counter[4] ;
 wire \simon1.tick_counter[5] ;
 wire \simon1.tick_counter[6] ;
 wire \simon1.tick_counter[7] ;
 wire \simon1.tick_counter[8] ;
 wire \simon1.tick_counter[9] ;
 wire \simon1.tone_sequence_counter[0] ;
 wire \simon1.tone_sequence_counter[1] ;
 wire \simon1.tone_sequence_counter[2] ;
 wire \simon1.user_input[0] ;
 wire \simon1.user_input[1] ;
 wire clknet_0_clk;
 wire net90;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_xnor2_1 _1313_ (.Y(_0247_),
    .A(_0244_),
    .B(_0246_));
 sg13g2_nor2_1 _1314_ (.A(net43),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_xnor2_1 _1315_ (.Y(_0249_),
    .A(\simon1.play1.tick_counter[4] ),
    .B(_0248_));
 sg13g2_nor2_1 _1316_ (.A(net77),
    .B(_0249_),
    .Y(_0102_));
 sg13g2_tiehi \simon1.millis_counter[8]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_xor2_1 _1318_ (.B(\simon1.play1.freq[5] ),
    .A(\simon1.play1.tick_counter[5] ),
    .X(_0251_));
 sg13g2_inv_1 _1319_ (.Y(_0252_),
    .A(\simon1.play1.freq[4] ));
 sg13g2_nor2_1 _1320_ (.A(_1043_),
    .B(_0240_),
    .Y(_0253_));
 sg13g2_nand2b_1 _1321_ (.Y(_0254_),
    .B(_0241_),
    .A_N(\simon1.play1.tick_counter[4] ));
 sg13g2_a22oi_1 _1322_ (.Y(_0255_),
    .B1(_0253_),
    .B2(_0254_),
    .A2(_0239_),
    .A1(_0237_));
 sg13g2_nor2_1 _1323_ (.A(\simon1.play1.tick_counter[4] ),
    .B(\simon1.play1.freq[4] ),
    .Y(_0256_));
 sg13g2_a22oi_1 _1324_ (.Y(_0257_),
    .B1(_0255_),
    .B2(_0256_),
    .A2(_0243_),
    .A1(_0252_));
 sg13g2_xor2_1 _1325_ (.B(_0257_),
    .A(_0251_),
    .X(_0258_));
 sg13g2_xor2_1 _1326_ (.B(_0232_),
    .A(\simon1.play1.freq[3] ),
    .X(_0259_));
 sg13g2_xor2_1 _1327_ (.B(\simon1.play1.freq[4] ),
    .A(\simon1.play1.tick_counter[4] ),
    .X(_0260_));
 sg13g2_and2_1 _1328_ (.A(\simon1.play1.tick_counter[3] ),
    .B(_0260_),
    .X(_0261_));
 sg13g2_nor4_1 _1329_ (.A(\simon1.play1.tick_counter[3] ),
    .B(net63),
    .C(_0232_),
    .D(_0260_),
    .Y(_0262_));
 sg13g2_and4_1 _1330_ (.A(_1043_),
    .B(net63),
    .C(_0232_),
    .D(_0260_),
    .X(_0263_));
 sg13g2_a22oi_1 _1331_ (.Y(_0264_),
    .B1(_0262_),
    .B2(_0263_),
    .A2(_0261_),
    .A1(_0259_));
 sg13g2_nand2_1 _1332_ (.Y(_0265_),
    .A(net34),
    .B(_0264_));
 sg13g2_xor2_1 _1333_ (.B(_0265_),
    .A(_0258_),
    .X(_0266_));
 sg13g2_nor2_1 _1334_ (.A(\simon1.play1.tick_counter[5] ),
    .B(net44),
    .Y(_0267_));
 sg13g2_tiehi \simon1.millis_counter[7]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_a22oi_1 _1336_ (.Y(_0103_),
    .B1(_0267_),
    .B2(net78),
    .A2(_0266_),
    .A1(net44));
 sg13g2_xnor2_1 _1337_ (.Y(_0269_),
    .A(\simon1.play1.tick_counter[6] ),
    .B(net62));
 sg13g2_a21o_1 _1338_ (.A2(_0239_),
    .A1(_0237_),
    .B1(_0242_),
    .X(_0270_));
 sg13g2_and2_1 _1339_ (.A(_0251_),
    .B(_0260_),
    .X(_0271_));
 sg13g2_nand2_1 _1340_ (.Y(_0272_),
    .A(\simon1.play1.tick_counter[4] ),
    .B(\simon1.play1.freq[4] ));
 sg13g2_nand2_1 _1341_ (.Y(_0273_),
    .A(\simon1.play1.tick_counter[5] ),
    .B(\simon1.play1.freq[5] ));
 sg13g2_nor2_1 _1342_ (.A(\simon1.play1.tick_counter[5] ),
    .B(\simon1.play1.freq[5] ),
    .Y(_0274_));
 sg13g2_a21oi_1 _1343_ (.A1(_0272_),
    .A2(_0273_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_a21oi_1 _1344_ (.A1(_0270_),
    .A2(_0271_),
    .Y(_0276_),
    .B1(_0275_));
 sg13g2_xor2_1 _1345_ (.B(_0276_),
    .A(_0269_),
    .X(_0277_));
 sg13g2_a21o_1 _1346_ (.A2(_0264_),
    .A1(_0258_),
    .B1(_1060_),
    .X(_0278_));
 sg13g2_xor2_1 _1347_ (.B(_0278_),
    .A(_0277_),
    .X(_0279_));
 sg13g2_nor2_1 _1348_ (.A(net43),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_a21oi_1 _1349_ (.A1(\simon1.play1.tick_counter[6] ),
    .A2(net43),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nor2_1 _1350_ (.A(net78),
    .B(_0281_),
    .Y(_0104_));
 sg13g2_xor2_1 _1351_ (.B(\simon1.play1.freq[7] ),
    .A(\simon1.play1.tick_counter[7] ),
    .X(_0282_));
 sg13g2_a21oi_1 _1352_ (.A1(\simon1.play1.tick_counter[6] ),
    .A2(net62),
    .Y(_0283_),
    .B1(_0282_));
 sg13g2_inv_1 _1353_ (.Y(_0284_),
    .A(_0282_));
 sg13g2_o21ai_1 _1354_ (.B1(\simon1.play1.tick_counter[6] ),
    .Y(_0285_),
    .A1(net62),
    .A2(_0275_));
 sg13g2_and2_1 _1355_ (.A(net62),
    .B(_0282_),
    .X(_0286_));
 sg13g2_nor2_1 _1356_ (.A(\simon1.play1.tick_counter[6] ),
    .B(net62),
    .Y(_0287_));
 sg13g2_nor2b_1 _1357_ (.A(_0282_),
    .B_N(_0287_),
    .Y(_0288_));
 sg13g2_a21oi_1 _1358_ (.A1(_0275_),
    .A2(_0286_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_o21ai_1 _1359_ (.B1(_0289_),
    .Y(_0290_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_inv_1 _1360_ (.Y(_0291_),
    .A(_0271_));
 sg13g2_nor4_1 _1361_ (.A(_0243_),
    .B(_0291_),
    .C(_0284_),
    .D(_0287_),
    .Y(_0292_));
 sg13g2_a22oi_1 _1362_ (.Y(_0293_),
    .B1(_0290_),
    .B2(_0292_),
    .A2(_0283_),
    .A1(_0276_));
 sg13g2_a21o_1 _1363_ (.A2(_0264_),
    .A1(_0258_),
    .B1(_0277_),
    .X(_0294_));
 sg13g2_tiehi \simon1.millis_counter[6]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_nand3_1 _1365_ (.B(_0293_),
    .C(_0294_),
    .A(net34),
    .Y(_0296_));
 sg13g2_a21o_1 _1366_ (.A2(_0294_),
    .A1(net34),
    .B1(_0293_),
    .X(_0297_));
 sg13g2_nand2_1 _1367_ (.Y(_0298_),
    .A(_0296_),
    .B(_0297_));
 sg13g2_nor2_1 _1368_ (.A(\simon1.play1.tick_counter[7] ),
    .B(_1075_),
    .Y(_0299_));
 sg13g2_a22oi_1 _1369_ (.Y(_0105_),
    .B1(_0299_),
    .B2(net78),
    .A2(_0298_),
    .A1(net45));
 sg13g2_xnor2_1 _1370_ (.Y(_0300_),
    .A(\simon1.play1.tick_counter[8] ),
    .B(\simon1.play1.freq[8] ));
 sg13g2_nor2b_1 _1371_ (.A(_0269_),
    .B_N(_0282_),
    .Y(_0301_));
 sg13g2_nand2_1 _1372_ (.Y(_0302_),
    .A(_0271_),
    .B(_0301_));
 sg13g2_nand3_1 _1373_ (.B(\simon1.play1.freq[5] ),
    .C(\simon1.play1.freq[6] ),
    .A(\simon1.play1.tick_counter[5] ),
    .Y(_0303_));
 sg13g2_a21oi_1 _1374_ (.A1(\simon1.play1.tick_counter[5] ),
    .A2(\simon1.play1.freq[5] ),
    .Y(_0304_),
    .B1(net62));
 sg13g2_nor2_1 _1375_ (.A(\simon1.play1.tick_counter[7] ),
    .B(\simon1.play1.freq[7] ),
    .Y(_0305_));
 sg13g2_a22oi_1 _1376_ (.Y(_0306_),
    .B1(_0304_),
    .B2(_0305_),
    .A2(_0303_),
    .A1(_1055_));
 sg13g2_and2_1 _1377_ (.A(\simon1.play1.tick_counter[7] ),
    .B(\simon1.play1.freq[7] ),
    .X(_0307_));
 sg13g2_nor4_1 _1378_ (.A(_0274_),
    .B(_0272_),
    .C(_0287_),
    .D(_0305_),
    .Y(_0308_));
 sg13g2_nor3_1 _1379_ (.A(_0306_),
    .B(_0307_),
    .C(_0308_),
    .Y(_0309_));
 sg13g2_o21ai_1 _1380_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_0243_),
    .A2(_0302_));
 sg13g2_xnor2_1 _1381_ (.Y(_0311_),
    .A(_0300_),
    .B(_0310_));
 sg13g2_xor2_1 _1382_ (.B(_0311_),
    .A(_0296_),
    .X(_0312_));
 sg13g2_nand3_1 _1383_ (.B(\simon1.play1.tick_counter[8] ),
    .C(net43),
    .A(net85),
    .Y(_0313_));
 sg13g2_o21ai_1 _1384_ (.B1(_0313_),
    .Y(_0106_),
    .A1(_1077_),
    .A2(_0312_));
 sg13g2_xor2_1 _1385_ (.B(\simon1.play1.freq[9] ),
    .A(\simon1.play1.tick_counter[9] ),
    .X(_0314_));
 sg13g2_o21ai_1 _1386_ (.B1(_0314_),
    .Y(_0315_),
    .A1(\simon1.play1.tick_counter[8] ),
    .A2(\simon1.play1.freq[8] ));
 sg13g2_nor3_1 _1387_ (.A(_0243_),
    .B(_0302_),
    .C(_0315_),
    .Y(_0316_));
 sg13g2_and2_1 _1388_ (.A(_0271_),
    .B(_0301_),
    .X(_0317_));
 sg13g2_or3_1 _1389_ (.A(_0306_),
    .B(_0307_),
    .C(_0308_),
    .X(_0318_));
 sg13g2_tiehi \simon1.millis_counter[5]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_and2_1 _1391_ (.A(\simon1.play1.tick_counter[8] ),
    .B(\simon1.play1.freq[8] ),
    .X(_0320_));
 sg13g2_or2_1 _1392_ (.X(_0321_),
    .B(_0320_),
    .A(_0314_));
 sg13g2_a22oi_1 _1393_ (.Y(_0322_),
    .B1(_0318_),
    .B2(_0321_),
    .A2(_0317_),
    .A1(_0270_));
 sg13g2_nor3_1 _1394_ (.A(\simon1.play1.tick_counter[8] ),
    .B(\simon1.play1.freq[8] ),
    .C(_0314_),
    .Y(_0323_));
 sg13g2_a21oi_1 _1395_ (.A1(_0314_),
    .A2(_0320_),
    .Y(_0324_),
    .B1(_0323_));
 sg13g2_o21ai_1 _1396_ (.B1(_0324_),
    .Y(_0325_),
    .A1(_0309_),
    .A2(_0315_));
 sg13g2_nor3_2 _1397_ (.A(_0316_),
    .B(_0322_),
    .C(_0325_),
    .Y(_0326_));
 sg13g2_and2_1 _1398_ (.A(_0293_),
    .B(_0311_),
    .X(_0327_));
 sg13g2_a21oi_1 _1399_ (.A1(_0294_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(net38));
 sg13g2_xnor2_1 _1400_ (.Y(_0329_),
    .A(_0326_),
    .B(_0328_));
 sg13g2_nor2_1 _1401_ (.A(\simon1.play1.tick_counter[9] ),
    .B(net44),
    .Y(_0330_));
 sg13g2_a22oi_1 _1402_ (.Y(_0107_),
    .B1(_0330_),
    .B2(net74),
    .A2(_0329_),
    .A1(net44));
 sg13g2_nand2b_2 _1403_ (.Y(_0331_),
    .B(_0314_),
    .A_N(_0300_));
 sg13g2_inv_1 _1404_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_a21oi_1 _1405_ (.A1(\simon1.play1.freq[9] ),
    .A2(_0320_),
    .Y(_0333_),
    .B1(\simon1.play1.tick_counter[9] ));
 sg13g2_nor2_1 _1406_ (.A(\simon1.play1.freq[9] ),
    .B(_0320_),
    .Y(_0334_));
 sg13g2_nor2_1 _1407_ (.A(_0333_),
    .B(_0334_),
    .Y(_0335_));
 sg13g2_a21o_2 _1408_ (.A2(_0332_),
    .A1(_0310_),
    .B1(_0335_),
    .X(_0336_));
 sg13g2_tiehi \simon1.millis_counter[4]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_nor2_1 _1410_ (.A(net42),
    .B(_0336_),
    .Y(_0338_));
 sg13g2_a22oi_1 _1411_ (.Y(_0339_),
    .B1(_0326_),
    .B2(net38),
    .A2(_0327_),
    .A1(_0294_));
 sg13g2_mux2_1 _1412_ (.A0(_0336_),
    .A1(_0338_),
    .S(_0339_),
    .X(_0340_));
 sg13g2_xnor2_1 _1413_ (.Y(_0341_),
    .A(\simon1.play1.tick_counter[10] ),
    .B(_0340_));
 sg13g2_nor2_1 _1414_ (.A(net74),
    .B(_0341_),
    .Y(_0108_));
 sg13g2_and2_1 _1415_ (.A(\simon1.play1.tick_counter[10] ),
    .B(_0336_),
    .X(_0342_));
 sg13g2_nor3_1 _1416_ (.A(\simon1.play1.tick_counter[10] ),
    .B(net42),
    .C(_0336_),
    .Y(_0343_));
 sg13g2_mux2_1 _1417_ (.A0(_0342_),
    .A1(_0343_),
    .S(_0339_),
    .X(_0344_));
 sg13g2_xnor2_1 _1418_ (.Y(_0345_),
    .A(\simon1.play1.tick_counter[11] ),
    .B(_0344_));
 sg13g2_nor2_1 _1419_ (.A(net78),
    .B(_0345_),
    .Y(_0109_));
 sg13g2_nand3b_1 _1420_ (.B(_0336_),
    .C(\simon1.play1.tick_counter[12] ),
    .Y(_0346_),
    .A_N(\simon1.play1.tick_counter[11] ));
 sg13g2_nand3_1 _1421_ (.B(\simon1.play1.tick_counter[10] ),
    .C(_0336_),
    .A(\simon1.play1.tick_counter[11] ),
    .Y(_0347_));
 sg13g2_mux2_1 _1422_ (.A0(_0347_),
    .A1(\simon1.play1.tick_counter[11] ),
    .S(\simon1.play1.tick_counter[12] ),
    .X(_0348_));
 sg13g2_a21o_1 _1423_ (.A2(_0346_),
    .A1(_0339_),
    .B1(_0348_),
    .X(_0349_));
 sg13g2_nand3_1 _1424_ (.B(\simon1.play1.tick_counter[11] ),
    .C(\simon1.play1.tick_counter[10] ),
    .A(\simon1.play1.tick_counter[12] ),
    .Y(_0350_));
 sg13g2_tiehi \simon1.millis_counter[3]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_nor4_1 _1426_ (.A(_0243_),
    .B(_0302_),
    .C(_0331_),
    .D(_0350_),
    .Y(_0352_));
 sg13g2_nor3_1 _1427_ (.A(_0309_),
    .B(_0331_),
    .C(_0350_),
    .Y(_0353_));
 sg13g2_nor3_1 _1428_ (.A(_0333_),
    .B(_0334_),
    .C(_0350_),
    .Y(_0354_));
 sg13g2_nor3_2 _1429_ (.A(_0352_),
    .B(_0353_),
    .C(_0354_),
    .Y(_0355_));
 sg13g2_a21oi_1 _1430_ (.A1(_0270_),
    .A2(_0317_),
    .Y(_0356_),
    .B1(_0318_));
 sg13g2_nor2_1 _1431_ (.A(_1037_),
    .B(_0335_),
    .Y(_0357_));
 sg13g2_o21ai_1 _1432_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0356_),
    .A2(_0331_));
 sg13g2_a221oi_1 _1433_ (.B2(_0358_),
    .C1(_0326_),
    .B1(_0355_),
    .A1(_0294_),
    .Y(_0359_),
    .A2(_0327_));
 sg13g2_tiehi \simon1.millis_counter[2]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_o21ai_1 _1435_ (.B1(\simon1.play1.tick_counter[12] ),
    .Y(_0361_),
    .A1(\simon1.play1.tick_counter[11] ),
    .A2(\simon1.play1.tick_counter[10] ));
 sg13g2_nor2b_1 _1436_ (.A(_0361_),
    .B_N(_0347_),
    .Y(_0362_));
 sg13g2_a22oi_1 _1437_ (.Y(_0363_),
    .B1(_0362_),
    .B2(net42),
    .A2(_0359_),
    .A1(net34));
 sg13g2_nor2_1 _1438_ (.A(\simon1.play1.tick_counter[12] ),
    .B(net44),
    .Y(_0364_));
 sg13g2_a22oi_1 _1439_ (.Y(_0110_),
    .B1(_0364_),
    .B2(net74),
    .A2(_0363_),
    .A1(_0349_));
 sg13g2_nor2_1 _1440_ (.A(net38),
    .B(_0359_),
    .Y(_0365_));
 sg13g2_or3_1 _1441_ (.A(_0352_),
    .B(_0353_),
    .C(_0354_),
    .X(_0366_));
 sg13g2_xnor2_1 _1442_ (.Y(_0367_),
    .A(_0034_),
    .B(_0366_));
 sg13g2_xnor2_1 _1443_ (.Y(_0368_),
    .A(_0365_),
    .B(_0367_));
 sg13g2_nor2_1 _1444_ (.A(\simon1.play1.tick_counter[13] ),
    .B(net45),
    .Y(_0369_));
 sg13g2_a22oi_1 _1445_ (.Y(_0111_),
    .B1(_0369_),
    .B2(net73),
    .A2(_0368_),
    .A1(net45));
 sg13g2_a21o_1 _1446_ (.A2(_0358_),
    .A1(_0355_),
    .B1(_0326_),
    .X(_0370_));
 sg13g2_a21o_1 _1447_ (.A2(_0327_),
    .A1(_0294_),
    .B1(_0370_),
    .X(_0371_));
 sg13g2_nor2_1 _1448_ (.A(\simon1.play1.tick_counter[13] ),
    .B(_0355_),
    .Y(_0372_));
 sg13g2_xnor2_1 _1449_ (.Y(_0373_),
    .A(_0034_),
    .B(_0372_));
 sg13g2_nand4_1 _1450_ (.B(net34),
    .C(_0371_),
    .A(net45),
    .Y(_0374_),
    .D(_0373_));
 sg13g2_inv_1 _1451_ (.Y(_0375_),
    .A(\simon1.play1.tick_counter[13] ));
 sg13g2_nor2_1 _1452_ (.A(_0375_),
    .B(_0355_),
    .Y(_0376_));
 sg13g2_o21ai_1 _1453_ (.B1(_0376_),
    .Y(_0377_),
    .A1(net38),
    .A2(_0359_));
 sg13g2_and3_1 _1454_ (.X(_0378_),
    .A(_1052_),
    .B(_0374_),
    .C(_0377_));
 sg13g2_a21oi_1 _1455_ (.A1(_0374_),
    .A2(_0377_),
    .Y(_0379_),
    .B1(_1052_));
 sg13g2_nor3_1 _1456_ (.A(net74),
    .B(_0378_),
    .C(_0379_),
    .Y(_0112_));
 sg13g2_nor2_1 _1457_ (.A(_1038_),
    .B(_0350_),
    .Y(_0380_));
 sg13g2_nand2_1 _1458_ (.Y(_0381_),
    .A(_0336_),
    .B(_0380_));
 sg13g2_nand2b_1 _1459_ (.Y(_0382_),
    .B(net81),
    .A_N(\simon1.play1.tick_counter[15] ));
 sg13g2_nor2_1 _1460_ (.A(_0381_),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_a22oi_1 _1461_ (.Y(_0384_),
    .B1(_0318_),
    .B2(_0335_),
    .A2(_0317_),
    .A1(_0270_));
 sg13g2_o21ai_1 _1462_ (.B1(_0380_),
    .Y(_0385_),
    .A1(_0335_),
    .A2(_0332_));
 sg13g2_nor2_2 _1463_ (.A(_0384_),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_nand2_1 _1464_ (.Y(_0387_),
    .A(net81),
    .B(\simon1.play1.tick_counter[15] ));
 sg13g2_nor2_1 _1465_ (.A(_0386_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_and4_1 _1466_ (.A(_1052_),
    .B(\simon1.play1.tick_counter[13] ),
    .C(_0034_),
    .D(_0366_),
    .X(_0389_));
 sg13g2_nand2b_1 _1467_ (.Y(_0390_),
    .B(\simon1.play1.tick_counter[14] ),
    .A_N(_0034_));
 sg13g2_nand3_1 _1468_ (.B(_0375_),
    .C(_0034_),
    .A(\simon1.play1.tick_counter[14] ),
    .Y(_0391_));
 sg13g2_mux2_1 _1469_ (.A0(_0390_),
    .A1(_0391_),
    .S(_0366_),
    .X(_0392_));
 sg13g2_nor2b_1 _1470_ (.A(_0389_),
    .B_N(_0392_),
    .Y(_0393_));
 sg13g2_o21ai_1 _1471_ (.B1(net34),
    .Y(_0394_),
    .A1(_0359_),
    .A2(_0393_));
 sg13g2_o21ai_1 _1472_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0383_),
    .A2(_0388_));
 sg13g2_a21oi_1 _1473_ (.A1(net44),
    .A2(_0381_),
    .Y(_0396_),
    .B1(_0387_));
 sg13g2_nand2b_1 _1474_ (.Y(_0397_),
    .B(_0396_),
    .A_N(_0394_));
 sg13g2_nand2_1 _1475_ (.Y(_0398_),
    .A(net44),
    .B(_0381_));
 sg13g2_or3_1 _1476_ (.A(_0394_),
    .B(_0398_),
    .C(_0382_),
    .X(_0399_));
 sg13g2_nand3_1 _1477_ (.B(_0397_),
    .C(_0399_),
    .A(_0395_),
    .Y(_0113_));
 sg13g2_nor2_1 _1478_ (.A(_0359_),
    .B(_0393_),
    .Y(_0400_));
 sg13g2_tiehi \simon1.millis_counter[1]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_or2_1 _1480_ (.X(_0402_),
    .B(\simon1.play1.tick_counter[16] ),
    .A(\simon1.play1.tick_counter[15] ));
 sg13g2_nor3_1 _1481_ (.A(net38),
    .B(_0398_),
    .C(_0402_),
    .Y(_0403_));
 sg13g2_nand2b_1 _1482_ (.Y(_0404_),
    .B(_0403_),
    .A_N(net22));
 sg13g2_or2_1 _1483_ (.X(_0405_),
    .B(_0398_),
    .A(\simon1.play1.tick_counter[15] ));
 sg13g2_o21ai_1 _1484_ (.B1(\simon1.play1.tick_counter[16] ),
    .Y(_0406_),
    .A1(_0400_),
    .A2(_0405_));
 sg13g2_a21oi_1 _1485_ (.A1(_0404_),
    .A2(_0406_),
    .Y(_0114_),
    .B1(net74));
 sg13g2_and2_1 _1486_ (.A(net81),
    .B(\simon1.play1.tick_counter[17] ),
    .X(_0407_));
 sg13g2_nor2_1 _1487_ (.A(net75),
    .B(\simon1.play1.tick_counter[17] ),
    .Y(_0408_));
 sg13g2_nor2b_1 _1488_ (.A(_0400_),
    .B_N(_0403_),
    .Y(_0409_));
 sg13g2_mux2_1 _1489_ (.A0(_0407_),
    .A1(_0408_),
    .S(_0409_),
    .X(_0115_));
 sg13g2_nand2_1 _1490_ (.Y(_0410_),
    .A(net81),
    .B(\simon1.play1.tick_counter[18] ));
 sg13g2_nor3_1 _1491_ (.A(\simon1.play1.tick_counter[17] ),
    .B(_0386_),
    .C(_0402_),
    .Y(_0411_));
 sg13g2_o21ai_1 _1492_ (.B1(_0411_),
    .Y(_0412_),
    .A1(_0359_),
    .A2(_0393_));
 sg13g2_nand4_1 _1493_ (.B(\simon1.play1.tick_counter[17] ),
    .C(\simon1.play1.tick_counter[16] ),
    .A(\simon1.play1.tick_counter[15] ),
    .Y(_0413_),
    .D(_0386_));
 sg13g2_a21oi_1 _1494_ (.A1(_0412_),
    .A2(_0413_),
    .Y(_0414_),
    .B1(net42));
 sg13g2_or3_1 _1495_ (.A(\simon1.play1.tick_counter[18] ),
    .B(\simon1.play1.tick_counter[17] ),
    .C(_0402_),
    .X(_0415_));
 sg13g2_nor2_1 _1496_ (.A(_0386_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nand2_1 _1497_ (.Y(_0417_),
    .A(net34),
    .B(_0416_));
 sg13g2_nand4_1 _1498_ (.B(\simon1.play1.tick_counter[18] ),
    .C(\simon1.play1.tick_counter[17] ),
    .A(\simon1.play1.tick_counter[15] ),
    .Y(_0418_),
    .D(\simon1.play1.tick_counter[16] ));
 sg13g2_or3_2 _1499_ (.A(_0384_),
    .B(_0385_),
    .C(_0418_),
    .X(_0419_));
 sg13g2_tiehi \simon1.millis_counter[0]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_a21oi_1 _1501_ (.A1(_0417_),
    .A2(_0419_),
    .Y(_0421_),
    .B1(_1077_));
 sg13g2_nand2b_1 _1502_ (.Y(_0422_),
    .B(_0421_),
    .A_N(net22));
 sg13g2_o21ai_1 _1503_ (.B1(_0422_),
    .Y(_0116_),
    .A1(_0410_),
    .A2(_0414_));
 sg13g2_nand2b_1 _1504_ (.Y(_0423_),
    .B(_0392_),
    .A_N(_0389_));
 sg13g2_a22oi_1 _1505_ (.Y(_0424_),
    .B1(_0417_),
    .B2(net42),
    .A2(_0423_),
    .A1(_0371_));
 sg13g2_tiehi _2444__101 (.L_HI(net101));
 sg13g2_xnor2_1 _1507_ (.Y(_0426_),
    .A(\simon1.play1.tick_counter[19] ),
    .B(net21));
 sg13g2_nor2_1 _1508_ (.A(net73),
    .B(_0426_),
    .Y(_0117_));
 sg13g2_nor4_1 _1509_ (.A(\simon1.play1.tick_counter[19] ),
    .B(net22),
    .C(_0398_),
    .D(_0415_),
    .Y(_0427_));
 sg13g2_nand2_1 _1510_ (.Y(_0428_),
    .A(net80),
    .B(\simon1.play1.tick_counter[20] ));
 sg13g2_nor2_1 _1511_ (.A(\simon1.play1.tick_counter[20] ),
    .B(\simon1.play1.tick_counter[19] ),
    .Y(_0429_));
 sg13g2_nand3_1 _1512_ (.B(_0429_),
    .C(net21),
    .A(net80),
    .Y(_0430_));
 sg13g2_o21ai_1 _1513_ (.B1(_0430_),
    .Y(_0118_),
    .A1(_0427_),
    .A2(_0428_));
 sg13g2_inv_1 _1514_ (.Y(_0431_),
    .A(\simon1.play1.tick_counter[21] ));
 sg13g2_a21o_1 _1515_ (.A2(net21),
    .A1(_0429_),
    .B1(_0431_),
    .X(_0432_));
 sg13g2_nand3_1 _1516_ (.B(_0429_),
    .C(net21),
    .A(_0431_),
    .Y(_0433_));
 sg13g2_a21oi_1 _1517_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0119_),
    .B1(net73));
 sg13g2_nor2_1 _1518_ (.A(net73),
    .B(\simon1.play1.tick_counter[22] ),
    .Y(_0434_));
 sg13g2_and2_1 _1519_ (.A(net80),
    .B(\simon1.play1.tick_counter[22] ),
    .X(_0435_));
 sg13g2_mux2_1 _1520_ (.A0(_0434_),
    .A1(_0435_),
    .S(_0433_),
    .X(_0120_));
 sg13g2_nand2_1 _1521_ (.Y(_0436_),
    .A(net80),
    .B(\simon1.play1.tick_counter[23] ));
 sg13g2_nor3_1 _1522_ (.A(_1025_),
    .B(_0386_),
    .C(_0415_),
    .Y(_0437_));
 sg13g2_o21ai_1 _1523_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0359_),
    .A2(_0393_));
 sg13g2_and4_1 _1524_ (.A(\simon1.play1.tick_counter[22] ),
    .B(\simon1.play1.tick_counter[21] ),
    .C(\simon1.play1.tick_counter[20] ),
    .D(\simon1.play1.tick_counter[19] ),
    .X(_0439_));
 sg13g2_nand2b_1 _1525_ (.Y(_0440_),
    .B(_0439_),
    .A_N(_0419_));
 sg13g2_a21oi_1 _1526_ (.A1(_0438_),
    .A2(_0440_),
    .Y(_0441_),
    .B1(net42));
 sg13g2_nor2_1 _1527_ (.A(_1026_),
    .B(net38),
    .Y(_0442_));
 sg13g2_nand2_1 _1528_ (.Y(_0443_),
    .A(\simon1.play1.tick_counter[23] ),
    .B(_0439_));
 sg13g2_nor2_1 _1529_ (.A(_0419_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_1 _1530_ (.A1(_0416_),
    .A2(_0442_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_or3_1 _1531_ (.A(_1077_),
    .B(net22),
    .C(_0445_),
    .X(_0446_));
 sg13g2_o21ai_1 _1532_ (.B1(_0446_),
    .Y(_0121_),
    .A1(_0436_),
    .A2(_0441_));
 sg13g2_nor2_1 _1533_ (.A(\simon1.play1.tick_counter[23] ),
    .B(_1025_),
    .Y(_0447_));
 sg13g2_inv_1 _1534_ (.Y(_0448_),
    .A(\simon1.play1.tick_counter[24] ));
 sg13g2_a21o_1 _1535_ (.A2(net21),
    .A1(_0447_),
    .B1(_0448_),
    .X(_0449_));
 sg13g2_nand3_1 _1536_ (.B(_0447_),
    .C(net21),
    .A(_0448_),
    .Y(_0450_));
 sg13g2_a21oi_1 _1537_ (.A1(_0449_),
    .A2(_0450_),
    .Y(_0122_),
    .B1(net73));
 sg13g2_nor2_1 _1538_ (.A(\simon1.play1.tick_counter[24] ),
    .B(_1026_),
    .Y(_0451_));
 sg13g2_inv_1 _1539_ (.Y(_0452_),
    .A(\simon1.play1.tick_counter[25] ));
 sg13g2_a21o_1 _1540_ (.A2(net21),
    .A1(_0451_),
    .B1(_0452_),
    .X(_0453_));
 sg13g2_nand3_1 _1541_ (.B(_0451_),
    .C(net21),
    .A(_0452_),
    .Y(_0454_));
 sg13g2_a21oi_1 _1542_ (.A1(_0453_),
    .A2(_0454_),
    .Y(_0123_),
    .B1(net73));
 sg13g2_nor4_2 _1543_ (.A(_0452_),
    .B(_0448_),
    .C(_0419_),
    .Y(_0455_),
    .D(_0443_));
 sg13g2_and2_1 _1544_ (.A(_1027_),
    .B(_0419_),
    .X(_0456_));
 sg13g2_a21oi_1 _1545_ (.A1(\simon1.play1.tick_counter[26] ),
    .A2(_0455_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_nand4_1 _1546_ (.B(net45),
    .C(_0451_),
    .A(_0452_),
    .Y(_0458_),
    .D(_0416_));
 sg13g2_inv_1 _1547_ (.Y(_0459_),
    .A(\simon1.play1.tick_counter[26] ));
 sg13g2_nor3_1 _1548_ (.A(net74),
    .B(_0459_),
    .C(_0455_),
    .Y(_0460_));
 sg13g2_o21ai_1 _1549_ (.B1(_0460_),
    .Y(_0461_),
    .A1(net22),
    .A2(_0458_));
 sg13g2_o21ai_1 _1550_ (.B1(_0461_),
    .Y(_0124_),
    .A1(_0422_),
    .A2(_0457_));
 sg13g2_nand2_1 _1551_ (.Y(_0462_),
    .A(_1027_),
    .B(_0416_));
 sg13g2_a22oi_1 _1552_ (.Y(_0463_),
    .B1(_0462_),
    .B2(net42),
    .A2(_0423_),
    .A1(_0371_));
 sg13g2_nand3b_1 _1553_ (.B(net34),
    .C(_0463_),
    .Y(_0464_),
    .A_N(\simon1.play1.tick_counter[27] ));
 sg13g2_nand2b_1 _1554_ (.Y(_0465_),
    .B(\simon1.play1.tick_counter[27] ),
    .A_N(_0463_));
 sg13g2_a21oi_1 _1555_ (.A1(_0464_),
    .A2(_0465_),
    .Y(_0125_),
    .B1(net74));
 sg13g2_nand3_1 _1556_ (.B(\simon1.play1.tick_counter[26] ),
    .C(_0455_),
    .A(\simon1.play1.tick_counter[27] ),
    .Y(_0466_));
 sg13g2_nand3_1 _1557_ (.B(\simon1.play1.tick_counter[28] ),
    .C(_0466_),
    .A(net80),
    .Y(_0467_));
 sg13g2_nor4_1 _1558_ (.A(\simon1.play1.tick_counter[27] ),
    .B(net42),
    .C(net22),
    .D(_0462_),
    .Y(_0468_));
 sg13g2_nor2_1 _1559_ (.A(\simon1.play1.tick_counter[28] ),
    .B(\simon1.play1.tick_counter[27] ),
    .Y(_0469_));
 sg13g2_and4_1 _1560_ (.A(\simon1.play1.tick_counter[28] ),
    .B(\simon1.play1.tick_counter[27] ),
    .C(\simon1.play1.tick_counter[26] ),
    .D(_0455_),
    .X(_0470_));
 sg13g2_a21o_1 _1561_ (.A2(_0456_),
    .A1(_0469_),
    .B1(_0470_),
    .X(_0471_));
 sg13g2_nand3b_1 _1562_ (.B(_0421_),
    .C(_0471_),
    .Y(_0472_),
    .A_N(net22));
 sg13g2_o21ai_1 _1563_ (.B1(_0472_),
    .Y(_0126_),
    .A1(_0467_),
    .A2(_0468_));
 sg13g2_and2_1 _1564_ (.A(net80),
    .B(\simon1.play1.tick_counter[29] ),
    .X(_0473_));
 sg13g2_nor2_1 _1565_ (.A(net73),
    .B(\simon1.play1.tick_counter[29] ),
    .Y(_0474_));
 sg13g2_nor2_1 _1566_ (.A(_0243_),
    .B(_0302_),
    .Y(_0475_));
 sg13g2_or2_1 _1567_ (.X(_0476_),
    .B(_0350_),
    .A(_1038_));
 sg13g2_nor3_1 _1568_ (.A(_0331_),
    .B(_0476_),
    .C(_0418_),
    .Y(_0477_));
 sg13g2_and2_1 _1569_ (.A(_0318_),
    .B(_0477_),
    .X(_0478_));
 sg13g2_nor4_1 _1570_ (.A(_0333_),
    .B(_0334_),
    .C(_0476_),
    .D(_0418_),
    .Y(_0479_));
 sg13g2_a22oi_1 _1571_ (.Y(_0480_),
    .B1(_0478_),
    .B2(_0479_),
    .A2(_0477_),
    .A1(_0475_));
 sg13g2_nand4_1 _1572_ (.B(_1027_),
    .C(_0469_),
    .A(net45),
    .Y(_0481_),
    .D(_0480_));
 sg13g2_a22oi_1 _1573_ (.Y(_0482_),
    .B1(_0481_),
    .B2(net22),
    .A2(_0419_),
    .A1(_0417_));
 sg13g2_mux2_1 _1574_ (.A0(_0473_),
    .A1(_0474_),
    .S(_0482_),
    .X(_0127_));
 sg13g2_and2_1 _1575_ (.A(\simon1.play1.tick_counter[30] ),
    .B(\simon1.play1.tick_counter[29] ),
    .X(_0483_));
 sg13g2_and2_1 _1576_ (.A(_1030_),
    .B(_0419_),
    .X(_0484_));
 sg13g2_a21oi_1 _1577_ (.A1(_0470_),
    .A2(_0483_),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_and4_1 _1578_ (.A(\simon1.play1.tick_counter[29] ),
    .B(\simon1.play1.tick_counter[28] ),
    .C(\simon1.play1.tick_counter[27] ),
    .D(\simon1.play1.tick_counter[26] ),
    .X(_0486_));
 sg13g2_nand3_1 _1579_ (.B(_0455_),
    .C(_0486_),
    .A(net45),
    .Y(_0487_));
 sg13g2_nand3_1 _1580_ (.B(\simon1.play1.tick_counter[30] ),
    .C(_0487_),
    .A(net80),
    .Y(_0488_));
 sg13g2_a21o_1 _1581_ (.A2(_0463_),
    .A1(_1029_),
    .B1(_0488_),
    .X(_0489_));
 sg13g2_o21ai_1 _1582_ (.B1(_0489_),
    .Y(_0128_),
    .A1(_0422_),
    .A2(_0485_));
 sg13g2_inv_1 _1583_ (.Y(_0490_),
    .A(\simon1.play1.tick_counter[31] ));
 sg13g2_a21o_1 _1584_ (.A2(_0424_),
    .A1(_1030_),
    .B1(_0490_),
    .X(_0491_));
 sg13g2_nand3_1 _1585_ (.B(_1030_),
    .C(_0424_),
    .A(_0490_),
    .Y(_0492_));
 sg13g2_a21oi_1 _1586_ (.A1(_0491_),
    .A2(_0492_),
    .Y(_0129_),
    .B1(net73));
 sg13g2_a21oi_1 _1587_ (.A1(\simon1.state[0] ),
    .A2(_0657_),
    .Y(_0493_),
    .B1(\simon1.score1.ena ));
 sg13g2_nor2_1 _1588_ (.A(net79),
    .B(_0493_),
    .Y(_0132_));
 sg13g2_and4_1 _1589_ (.A(net83),
    .B(_1124_),
    .C(net39),
    .D(net35),
    .X(_0133_));
 sg13g2_and2_1 _1590_ (.A(net81),
    .B(_0037_),
    .X(_0136_));
 sg13g2_xnor2_1 _1591_ (.Y(_0494_),
    .A(\simon1.next_random[0] ),
    .B(\simon1.next_random[1] ));
 sg13g2_nor2_1 _1592_ (.A(net75),
    .B(_0494_),
    .Y(_0137_));
 sg13g2_a21oi_1 _1593_ (.A1(_0033_),
    .A2(net40),
    .Y(_0495_),
    .B1(_0966_));
 sg13g2_nor2_1 _1594_ (.A(net49),
    .B(net40),
    .Y(_0496_));
 sg13g2_nor2_1 _1595_ (.A(_0963_),
    .B(_0657_),
    .Y(_0497_));
 sg13g2_o21ai_1 _1596_ (.B1(_0497_),
    .Y(_0498_),
    .A1(_0495_),
    .A2(_0496_));
 sg13g2_nor4_2 _1597_ (.A(\simon1.state[6] ),
    .B(\simon1.state[3] ),
    .C(net56),
    .Y(_0499_),
    .D(\simon1.state[7] ));
 sg13g2_nand2b_1 _1598_ (.Y(_0500_),
    .B(_0499_),
    .A_N(\simon1.state[2] ));
 sg13g2_nand2_1 _1599_ (.Y(_0501_),
    .A(net54),
    .B(_0814_));
 sg13g2_and4_2 _1600_ (.A(_0977_),
    .B(_0498_),
    .C(_0500_),
    .D(_0501_),
    .X(_0502_));
 sg13g2_tiehi _2443__100 (.L_HI(net100));
 sg13g2_xnor2_1 _1602_ (.Y(_0504_),
    .A(net51),
    .B(net48));
 sg13g2_nand3b_1 _1603_ (.B(net47),
    .C(net51),
    .Y(_0505_),
    .A_N(net48));
 sg13g2_o21ai_1 _1604_ (.B1(_0505_),
    .Y(_0506_),
    .A1(net53),
    .A2(_0504_));
 sg13g2_nand2_1 _1605_ (.Y(_0507_),
    .A(_0497_),
    .B(_0970_));
 sg13g2_nor2_1 _1606_ (.A(net64),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_a221oi_1 _1607_ (.B2(net58),
    .C1(_0508_),
    .B1(_0506_),
    .A1(net53),
    .Y(_0509_),
    .A2(_0497_));
 sg13g2_nor2_1 _1608_ (.A(\simon1.play1.freq[0] ),
    .B(_0502_),
    .Y(_0510_));
 sg13g2_a22oi_1 _1609_ (.Y(_0141_),
    .B1(_0510_),
    .B2(net77),
    .A2(_0509_),
    .A1(_0502_));
 sg13g2_inv_1 _1610_ (.Y(_0511_),
    .A(\simon1.play1.freq[1] ));
 sg13g2_nand4_1 _1611_ (.B(_0498_),
    .C(_0500_),
    .A(_0977_),
    .Y(_0512_),
    .D(_0501_));
 sg13g2_tiehi _2442__99 (.L_HI(net99));
 sg13g2_xor2_1 _1613_ (.B(net41),
    .A(_0706_),
    .X(_0514_));
 sg13g2_xnor2_1 _1614_ (.Y(_0515_),
    .A(\simon1.millis_counter[1] ),
    .B(net64));
 sg13g2_nand2_1 _1615_ (.Y(_0516_),
    .A(net49),
    .B(_0966_));
 sg13g2_a21oi_1 _1616_ (.A1(_0969_),
    .A2(_0515_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_xor2_1 _1617_ (.B(\simon1.user_input[1] ),
    .A(\simon1.user_input[0] ),
    .X(_0518_));
 sg13g2_nor2_1 _1618_ (.A(_0983_),
    .B(net50),
    .Y(_0519_));
 sg13g2_a22oi_1 _1619_ (.Y(_0520_),
    .B1(_0519_),
    .B2(_0873_),
    .A2(net48),
    .A1(net51));
 sg13g2_a21oi_1 _1620_ (.A1(_0772_),
    .A2(_0518_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_o21ai_1 _1621_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0663_),
    .A2(_0517_));
 sg13g2_a22oi_1 _1622_ (.Y(_0523_),
    .B1(_0522_),
    .B2(_0512_),
    .A2(_0514_),
    .A1(_0499_));
 sg13g2_a22oi_1 _1623_ (.Y(_0142_),
    .B1(_0523_),
    .B2(net77),
    .A2(_0512_),
    .A1(_0511_));
 sg13g2_o21ai_1 _1624_ (.B1(\simon1.millis_counter[2] ),
    .Y(_0524_),
    .A1(\simon1.millis_counter[1] ),
    .A2(\simon1.millis_counter[0] ));
 sg13g2_nand2_1 _1625_ (.Y(_0525_),
    .A(_0967_),
    .B(_0524_));
 sg13g2_a21oi_1 _1626_ (.A1(net49),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0663_));
 sg13g2_nor3_1 _1627_ (.A(_0771_),
    .B(\simon1.user_input[1] ),
    .C(net40),
    .Y(_0527_));
 sg13g2_a22oi_1 _1628_ (.Y(_0528_),
    .B1(_0527_),
    .B2(_0499_),
    .A2(_0526_),
    .A1(_0966_));
 sg13g2_and2_1 _1629_ (.A(_0706_),
    .B(_0499_),
    .X(_0529_));
 sg13g2_nor3_1 _1630_ (.A(net33),
    .B(_0528_),
    .C(_0529_),
    .Y(_0530_));
 sg13g2_a21oi_1 _1631_ (.A1(\simon1.play1.freq[2] ),
    .A2(net33),
    .Y(_0531_),
    .B1(_0530_));
 sg13g2_nor2_1 _1632_ (.A(net77),
    .B(_0531_),
    .Y(_0143_));
 sg13g2_nand2b_1 _1633_ (.Y(_0532_),
    .B(_0529_),
    .A_N(net41));
 sg13g2_nor2b_1 _1634_ (.A(\simon1.user_input[0] ),
    .B_N(\simon1.user_input[1] ),
    .Y(_0533_));
 sg13g2_nor2b_1 _1635_ (.A(net52),
    .B_N(net51),
    .Y(_0534_));
 sg13g2_a22oi_1 _1636_ (.Y(_0535_),
    .B1(_0534_),
    .B2(_0873_),
    .A2(net48),
    .A1(net53));
 sg13g2_xnor2_1 _1637_ (.Y(_0536_),
    .A(\simon1.millis_counter[3] ),
    .B(_0524_));
 sg13g2_a21oi_1 _1638_ (.A1(_0974_),
    .A2(_0536_),
    .Y(_0537_),
    .B1(_0663_));
 sg13g2_a22oi_1 _1639_ (.Y(_0538_),
    .B1(_0535_),
    .B2(_0537_),
    .A2(_0533_),
    .A1(_0772_));
 sg13g2_nand3_1 _1640_ (.B(_0532_),
    .C(_0538_),
    .A(_0502_),
    .Y(_0539_));
 sg13g2_o21ai_1 _1641_ (.B1(_0539_),
    .Y(_0540_),
    .A1(net63),
    .A2(_0502_));
 sg13g2_nor2_1 _1642_ (.A(net77),
    .B(_0540_),
    .Y(_0144_));
 sg13g2_and2_1 _1643_ (.A(\simon1.user_input[0] ),
    .B(\simon1.user_input[1] ),
    .X(_0541_));
 sg13g2_a221oi_1 _1644_ (.B2(_0772_),
    .C1(net33),
    .B1(_0541_),
    .A1(net41),
    .Y(_0542_),
    .A2(_0529_));
 sg13g2_mux2_1 _1645_ (.A0(_0534_),
    .A1(_0519_),
    .S(net48),
    .X(_0543_));
 sg13g2_nor2b_1 _1646_ (.A(\simon1.millis_counter[3] ),
    .B_N(_0524_),
    .Y(_0544_));
 sg13g2_xnor2_1 _1647_ (.Y(_0545_),
    .A(\simon1.millis_counter[4] ),
    .B(_0544_));
 sg13g2_nor2_1 _1648_ (.A(_0507_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_a21oi_1 _1649_ (.A1(net58),
    .A2(_0543_),
    .Y(_0547_),
    .B1(_0546_));
 sg13g2_a221oi_1 _1650_ (.B2(_0547_),
    .C1(net77),
    .B1(_0542_),
    .A1(_0252_),
    .Y(_0145_),
    .A2(net33));
 sg13g2_nand2_1 _1651_ (.Y(_0548_),
    .A(_0020_),
    .B(_0544_));
 sg13g2_a21o_1 _1652_ (.A2(_0548_),
    .A1(_0974_),
    .B1(_0499_),
    .X(_0549_));
 sg13g2_nor4_1 _1653_ (.A(net53),
    .B(_0035_),
    .C(_0657_),
    .D(_0549_),
    .Y(_0550_));
 sg13g2_mux2_1 _1654_ (.A0(\simon1.play1.freq[5] ),
    .A1(_0550_),
    .S(_0502_),
    .X(_0551_));
 sg13g2_and2_1 _1655_ (.A(net85),
    .B(_0551_),
    .X(_0146_));
 sg13g2_inv_1 _1656_ (.Y(_0552_),
    .A(net62));
 sg13g2_or4_1 _1657_ (.A(\simon1.state[6] ),
    .B(\simon1.state[3] ),
    .C(net56),
    .D(\simon1.state[7] ),
    .X(_0553_));
 sg13g2_nor2_1 _1658_ (.A(net41),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_a21oi_1 _1659_ (.A1(net47),
    .A2(net48),
    .Y(_0555_),
    .B1(_0966_));
 sg13g2_nand2b_1 _1660_ (.Y(_0556_),
    .B(_0772_),
    .A_N(\simon1.user_input[0] ));
 sg13g2_o21ai_1 _1661_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0873_),
    .A2(_0555_));
 sg13g2_nor3_1 _1662_ (.A(net51),
    .B(_0663_),
    .C(_0549_),
    .Y(_0558_));
 sg13g2_nor4_1 _1663_ (.A(net33),
    .B(_0554_),
    .C(_0557_),
    .D(_0558_),
    .Y(_0559_));
 sg13g2_a22oi_1 _1664_ (.Y(_0147_),
    .B1(_0559_),
    .B2(net78),
    .A2(net33),
    .A1(_0552_));
 sg13g2_o21ai_1 _1665_ (.B1(_0499_),
    .Y(_0560_),
    .A1(_0706_),
    .A2(net41));
 sg13g2_nor2_1 _1666_ (.A(_0873_),
    .B(net48),
    .Y(_0561_));
 sg13g2_o21ai_1 _1667_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0519_),
    .A2(_0534_));
 sg13g2_nor2_1 _1668_ (.A(\simon1.user_input[0] ),
    .B(\simon1.user_input[1] ),
    .Y(_0563_));
 sg13g2_nor2_1 _1669_ (.A(_0507_),
    .B(_0548_),
    .Y(_0564_));
 sg13g2_a21oi_1 _1670_ (.A1(_0772_),
    .A2(_0563_),
    .Y(_0565_),
    .B1(_0564_));
 sg13g2_nand3_1 _1671_ (.B(_0562_),
    .C(_0565_),
    .A(_0553_),
    .Y(_0566_));
 sg13g2_nand3_1 _1672_ (.B(_0560_),
    .C(_0566_),
    .A(_0502_),
    .Y(_0567_));
 sg13g2_nand2_1 _1673_ (.Y(_0568_),
    .A(\simon1.play1.freq[7] ),
    .B(net33));
 sg13g2_a21oi_1 _1674_ (.A1(_0567_),
    .A2(_0568_),
    .Y(_0148_),
    .B1(net78));
 sg13g2_nor3_1 _1675_ (.A(_0771_),
    .B(_0749_),
    .C(_0563_),
    .Y(_0569_));
 sg13g2_o21ai_1 _1676_ (.B1(net49),
    .Y(_0570_),
    .A1(_0983_),
    .A2(net47));
 sg13g2_a221oi_1 _1677_ (.B2(net50),
    .C1(_0873_),
    .B1(_0570_),
    .A1(net49),
    .Y(_0571_),
    .A2(_0026_));
 sg13g2_nor4_1 _1678_ (.A(net33),
    .B(_0564_),
    .C(_0569_),
    .D(_0571_),
    .Y(_0572_));
 sg13g2_o21ai_1 _1679_ (.B1(net85),
    .Y(_0573_),
    .A1(\simon1.play1.freq[8] ),
    .A2(_0502_));
 sg13g2_a21oi_1 _1680_ (.A1(_0560_),
    .A2(_0572_),
    .Y(_0149_),
    .B1(_0573_));
 sg13g2_a21o_1 _1681_ (.A2(_0548_),
    .A1(_0969_),
    .B1(_0516_),
    .X(_0574_));
 sg13g2_nor2_1 _1682_ (.A(_0873_),
    .B(_0504_),
    .Y(_0575_));
 sg13g2_a21oi_1 _1683_ (.A1(_0497_),
    .A2(_0574_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_o21ai_1 _1684_ (.B1(net85),
    .Y(_0577_),
    .A1(\simon1.play1.freq[9] ),
    .A2(_0502_));
 sg13g2_a21oi_1 _1685_ (.A1(_0542_),
    .A2(_0576_),
    .Y(_0150_),
    .B1(_0577_));
 sg13g2_a21oi_1 _1686_ (.A1(net55),
    .A2(_0739_),
    .Y(_0578_),
    .B1(net54));
 sg13g2_o21ai_1 _1687_ (.B1(_0977_),
    .Y(_0579_),
    .A1(_0771_),
    .A2(net40));
 sg13g2_nor3_1 _1688_ (.A(\simon1.state[0] ),
    .B(\simon1.state[1] ),
    .C(_0500_),
    .Y(_0580_));
 sg13g2_o21ai_1 _1689_ (.B1(\simon1.state[7] ),
    .Y(_0581_),
    .A1(_0814_),
    .A2(_0974_));
 sg13g2_a21oi_1 _1690_ (.A1(_0654_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(_0657_));
 sg13g2_nor4_1 _1691_ (.A(_0763_),
    .B(_0579_),
    .C(_0580_),
    .D(_0582_),
    .Y(_0583_));
 sg13g2_o21ai_1 _1692_ (.B1(_0583_),
    .Y(_0584_),
    .A1(_0812_),
    .A2(_0578_));
 sg13g2_nand2_1 _1693_ (.Y(_0585_),
    .A(net83),
    .B(_0584_));
 sg13g2_xnor2_1 _1694_ (.Y(_0586_),
    .A(net64),
    .B(_1084_));
 sg13g2_nor2_1 _1695_ (.A(_0585_),
    .B(_0586_),
    .Y(_0151_));
 sg13g2_and2_1 _1696_ (.A(_1084_),
    .B(_0515_),
    .X(_0587_));
 sg13g2_a22oi_1 _1697_ (.Y(_0152_),
    .B1(_0585_),
    .B2(_0587_),
    .A2(_1086_),
    .A1(_0017_));
 sg13g2_and2_2 _1698_ (.A(net83),
    .B(_0584_),
    .X(_0588_));
 sg13g2_tiehi _2441__98 (.L_HI(net98));
 sg13g2_nand3_1 _1700_ (.B(net64),
    .C(_1084_),
    .A(\simon1.millis_counter[1] ),
    .Y(_0590_));
 sg13g2_xor2_1 _1701_ (.B(_0590_),
    .A(_0018_),
    .X(_0591_));
 sg13g2_and2_1 _1702_ (.A(_0588_),
    .B(_0591_),
    .X(_0153_));
 sg13g2_nor2_1 _1703_ (.A(_0018_),
    .B(_0590_),
    .Y(_0592_));
 sg13g2_xnor2_1 _1704_ (.Y(_0593_),
    .A(_0019_),
    .B(_0592_));
 sg13g2_and2_1 _1705_ (.A(_0588_),
    .B(_0593_),
    .X(_0154_));
 sg13g2_nand4_1 _1706_ (.B(net64),
    .C(\simon1.millis_counter[3] ),
    .A(\simon1.millis_counter[1] ),
    .Y(_0594_),
    .D(\simon1.millis_counter[2] ));
 sg13g2_xnor2_1 _1707_ (.Y(_0595_),
    .A(\simon1.millis_counter[4] ),
    .B(_0594_));
 sg13g2_nor2_1 _1708_ (.A(_0020_),
    .B(_1084_),
    .Y(_0596_));
 sg13g2_a21oi_1 _1709_ (.A1(_1084_),
    .A2(_0595_),
    .Y(_0597_),
    .B1(_0596_));
 sg13g2_nor2b_1 _1710_ (.A(_0597_),
    .B_N(_0588_),
    .Y(_0155_));
 sg13g2_nor2_1 _1711_ (.A(_1086_),
    .B(_0594_),
    .Y(_0598_));
 sg13g2_nand2_1 _1712_ (.Y(_0599_),
    .A(\simon1.millis_counter[4] ),
    .B(_0598_));
 sg13g2_xor2_1 _1713_ (.B(_0599_),
    .A(_0021_),
    .X(_0600_));
 sg13g2_and2_1 _1714_ (.A(_0588_),
    .B(_0600_),
    .X(_0156_));
 sg13g2_nand2b_1 _1715_ (.Y(_0601_),
    .B(_0598_),
    .A_N(_0775_));
 sg13g2_xor2_1 _1716_ (.B(_0601_),
    .A(_0022_),
    .X(_0602_));
 sg13g2_and2_1 _1717_ (.A(_0588_),
    .B(_0602_),
    .X(_0157_));
 sg13g2_nor2_1 _1718_ (.A(_0022_),
    .B(_0601_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1719_ (.Y(_0604_),
    .A(_0023_),
    .B(_0603_));
 sg13g2_and2_1 _1720_ (.A(_0588_),
    .B(_0604_),
    .X(_0158_));
 sg13g2_or2_1 _1721_ (.X(_0605_),
    .B(_0601_),
    .A(_0774_));
 sg13g2_xor2_1 _1722_ (.B(_0605_),
    .A(_0024_),
    .X(_0606_));
 sg13g2_and2_1 _1723_ (.A(_0588_),
    .B(_0606_),
    .X(_0159_));
 sg13g2_nor2_1 _1724_ (.A(_0024_),
    .B(_0605_),
    .Y(_0607_));
 sg13g2_xnor2_1 _1725_ (.Y(_0608_),
    .A(_0025_),
    .B(_0607_));
 sg13g2_and2_1 _1726_ (.A(_0588_),
    .B(_0608_),
    .X(_0160_));
 sg13g2_nand2_1 _1727_ (.Y(_0609_),
    .A(_1124_),
    .B(_1128_));
 sg13g2_nand3_1 _1728_ (.B(net35),
    .C(_0609_),
    .A(net60),
    .Y(_0610_));
 sg13g2_o21ai_1 _1729_ (.B1(_0610_),
    .Y(_0611_),
    .A1(net60),
    .A2(net35));
 sg13g2_nor2_1 _1730_ (.A(_0032_),
    .B(net39),
    .Y(_0612_));
 sg13g2_a21oi_1 _1731_ (.A1(net35),
    .A2(_0612_),
    .Y(_0613_),
    .B1(_0874_));
 sg13g2_nor2_1 _1732_ (.A(net60),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_a22oi_1 _1733_ (.Y(_0177_),
    .B1(_0614_),
    .B2(net76),
    .A2(_0611_),
    .A1(net55));
 sg13g2_a21oi_1 _1734_ (.A1(net60),
    .A2(net35),
    .Y(_0615_),
    .B1(_0771_));
 sg13g2_o21ai_1 _1735_ (.B1(\simon1.seq_length[1] ),
    .Y(_0616_),
    .A1(_0874_),
    .A2(_0615_));
 sg13g2_nand2_1 _1736_ (.Y(_0617_),
    .A(net60),
    .B(net55));
 sg13g2_nor3_1 _1737_ (.A(\simon1.seq_length[1] ),
    .B(_0612_),
    .C(_0617_),
    .Y(_0618_));
 sg13g2_and2_1 _1738_ (.A(\simon1.seq_length[1] ),
    .B(_0612_),
    .X(_0619_));
 sg13g2_o21ai_1 _1739_ (.B1(net35),
    .Y(_0620_),
    .A1(_0618_),
    .A2(_0619_));
 sg13g2_a21oi_1 _1740_ (.A1(_0616_),
    .A2(_0620_),
    .Y(_0178_),
    .B1(net76));
 sg13g2_nand2_1 _1741_ (.Y(_0621_),
    .A(net60),
    .B(\simon1.seq_length[1] ));
 sg13g2_xnor2_1 _1742_ (.Y(_0622_),
    .A(_0029_),
    .B(_0621_));
 sg13g2_nand4_1 _1743_ (.B(net55),
    .C(net35),
    .A(net83),
    .Y(_0623_),
    .D(_0609_));
 sg13g2_a21oi_1 _1744_ (.A1(_1123_),
    .A2(_0613_),
    .Y(_0624_),
    .B1(net76));
 sg13g2_nand2_1 _1745_ (.Y(_0625_),
    .A(\simon1.seq_length[2] ),
    .B(_0624_));
 sg13g2_o21ai_1 _1746_ (.B1(_0625_),
    .Y(_0179_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_nor2_1 _1747_ (.A(_0029_),
    .B(_0621_),
    .Y(_0626_));
 sg13g2_xor2_1 _1748_ (.B(_0626_),
    .A(_0030_),
    .X(_0627_));
 sg13g2_nand2_1 _1749_ (.Y(_0628_),
    .A(\simon1.seq_length[3] ),
    .B(_0624_));
 sg13g2_o21ai_1 _1750_ (.B1(_0628_),
    .Y(_0180_),
    .A1(_0623_),
    .A2(_0627_));
 sg13g2_nor2_1 _1751_ (.A(_0900_),
    .B(_0621_),
    .Y(_0629_));
 sg13g2_xor2_1 _1752_ (.B(_0629_),
    .A(_0031_),
    .X(_0630_));
 sg13g2_nand2_1 _1753_ (.Y(_0631_),
    .A(\simon1.seq_length[4] ),
    .B(_0624_));
 sg13g2_o21ai_1 _1754_ (.B1(_0631_),
    .Y(_0181_),
    .A1(_0623_),
    .A2(_0630_));
 sg13g2_a21oi_2 _1755_ (.B1(\simon1.state[4] ),
    .Y(_0632_),
    .A2(_0814_),
    .A1(net54));
 sg13g2_o21ai_1 _1756_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_0758_),
    .A2(_0663_));
 sg13g2_nand3b_1 _1757_ (.B(_0823_),
    .C(_0662_),
    .Y(_0634_),
    .A_N(_0500_));
 sg13g2_nor2_1 _1758_ (.A(_0780_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_a22oi_1 _1759_ (.Y(_0636_),
    .B1(_0633_),
    .B2(_0635_),
    .A2(_0563_),
    .A1(net57));
 sg13g2_nand2b_1 _1760_ (.Y(_0637_),
    .B(\simon1.state[2] ),
    .A_N(net57));
 sg13g2_nor2_1 _1761_ (.A(_0706_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nand2b_1 _1762_ (.Y(_0639_),
    .B(_0638_),
    .A_N(_0736_));
 sg13g2_nor2_1 _1763_ (.A(net14),
    .B(_0632_),
    .Y(_0640_));
 sg13g2_a22oi_1 _1764_ (.Y(_0182_),
    .B1(_0640_),
    .B2(net79),
    .A2(_0639_),
    .A1(_0636_));
 sg13g2_nand3b_1 _1765_ (.B(\simon1.user_input[0] ),
    .C(net57),
    .Y(_0641_),
    .A_N(\simon1.user_input[1] ));
 sg13g2_o21ai_1 _1766_ (.B1(_0641_),
    .Y(_0642_),
    .A1(_0744_),
    .A2(_0634_));
 sg13g2_a22oi_1 _1767_ (.Y(_0643_),
    .B1(_0642_),
    .B2(_0633_),
    .A2(_0638_),
    .A1(_0736_));
 sg13g2_o21ai_1 _1768_ (.B1(net85),
    .Y(_0644_),
    .A1(net15),
    .A2(_0632_));
 sg13g2_nor2_1 _1769_ (.A(_0643_),
    .B(_0644_),
    .Y(_0183_));
 sg13g2_o21ai_1 _1770_ (.B1(net85),
    .Y(_0645_),
    .A1(net16),
    .A2(_0632_));
 sg13g2_nand2b_1 _1771_ (.Y(_0646_),
    .B(_0706_),
    .A_N(_0637_));
 sg13g2_a21oi_1 _1772_ (.A1(\simon1.millis_counter[9] ),
    .A2(_0743_),
    .Y(_0647_),
    .B1(_0634_));
 sg13g2_a22oi_1 _1773_ (.Y(_0648_),
    .B1(_0633_),
    .B2(_0647_),
    .A2(_0533_),
    .A1(net57));
 sg13g2_o21ai_1 _1774_ (.B1(_0648_),
    .Y(_0649_),
    .A1(net41),
    .A2(_0646_));
 sg13g2_nor2b_1 _1775_ (.A(_0645_),
    .B_N(_0649_),
    .Y(_0184_));
 sg13g2_nor2b_1 _1776_ (.A(_0634_),
    .B_N(_0968_),
    .Y(_0650_));
 sg13g2_a22oi_1 _1777_ (.Y(_0651_),
    .B1(_0633_),
    .B2(_0650_),
    .A2(_0541_),
    .A1(net57));
 sg13g2_nand2b_1 _1778_ (.Y(_0652_),
    .B(net41),
    .A_N(_0646_));
 sg13g2_nor2_1 _1779_ (.A(net17),
    .B(_0632_),
    .Y(_0653_));
 sg13g2_a22oi_1 _1780_ (.Y(_0185_),
    .B1(_0653_),
    .B2(net76),
    .A2(_0652_),
    .A1(_0651_));
 sg13g2_inv_1 _1781_ (.Y(_0654_),
    .A(\simon1.state[0] ));
 sg13g2_nor2_1 _1782_ (.A(net4),
    .B(net5),
    .Y(_0655_));
 sg13g2_nor2_1 _1783_ (.A(net2),
    .B(net3),
    .Y(_0656_));
 sg13g2_nand2_2 _1784_ (.Y(_0657_),
    .A(_0655_),
    .B(_0656_));
 sg13g2_tiehi _2440__97 (.L_HI(net97));
 sg13g2_tiehi _2439__96 (.L_HI(net96));
 sg13g2_tiehi _2435__95 (.L_HI(net95));
 sg13g2_o21ai_1 _1788_ (.B1(net83),
    .Y(_0005_),
    .A1(_0654_),
    .A2(_0657_));
 sg13g2_tiehi _2434__94 (.L_HI(net94));
 sg13g2_and2_1 _1790_ (.A(_0655_),
    .B(_0656_),
    .X(_0662_));
 sg13g2_nand2_2 _1791_ (.Y(_0663_),
    .A(\simon1.state[7] ),
    .B(_0662_));
 sg13g2_tiehi _2433__93 (.L_HI(net93));
 sg13g2_tiehi _2432__92 (.L_HI(net92));
 sg13g2_tiehi _2431__91 (.L_HI(net91));
 sg13g2_tielo _2448__89 (.L_LO(net89));
 sg13g2_tielo _2446__88 (.L_LO(net88));
 sg13g2_mux4_1 _1797_ (.S0(net71),
    .A0(\simon1.seq[12][1] ),
    .A1(\simon1.seq[13][1] ),
    .A2(\simon1.seq[14][1] ),
    .A3(\simon1.seq[15][1] ),
    .S1(net68),
    .X(_0669_));
 sg13g2_mux4_1 _1798_ (.S0(net72),
    .A0(\simon1.seq[28][1] ),
    .A1(\simon1.seq[29][1] ),
    .A2(\simon1.seq[30][1] ),
    .A3(\simon1.seq[31][1] ),
    .S1(net70),
    .X(_0670_));
 sg13g2_tielo ttsimon_87 (.L_LO(net87));
 sg13g2_mux2_1 _1800_ (.A0(_0669_),
    .A1(_0670_),
    .S(_0004_),
    .X(_0672_));
 sg13g2_nand3_1 _1801_ (.B(_0003_),
    .C(_0672_),
    .A(_0002_),
    .Y(_0673_));
 sg13g2_nor2b_1 _1802_ (.A(_0002_),
    .B_N(_0003_),
    .Y(_0674_));
 sg13g2_buf_1 fanout86 (.A(net1),
    .X(net86));
 sg13g2_mux4_1 _1804_ (.S0(net71),
    .A0(\simon1.seq[8][1] ),
    .A1(\simon1.seq[9][1] ),
    .A2(\simon1.seq[10][1] ),
    .A3(\simon1.seq[11][1] ),
    .S1(net68),
    .X(_0676_));
 sg13g2_mux4_1 _1805_ (.S0(net71),
    .A0(\simon1.seq[24][1] ),
    .A1(\simon1.seq[25][1] ),
    .A2(\simon1.seq[26][1] ),
    .A3(\simon1.seq[27][1] ),
    .S1(net68),
    .X(_0677_));
 sg13g2_mux2_1 _1806_ (.A0(_0676_),
    .A1(_0677_),
    .S(_0004_),
    .X(_0678_));
 sg13g2_nand2_1 _1807_ (.Y(_0679_),
    .A(_0674_),
    .B(_0678_));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_nand2_2 _1809_ (.Y(_0681_),
    .A(net72),
    .B(_0004_));
 sg13g2_nor2b_1 _1810_ (.A(net66),
    .B_N(\simon1.seq[17][1] ),
    .Y(_0682_));
 sg13g2_a22oi_1 _1811_ (.Y(_0683_),
    .B1(_0681_),
    .B2(_0682_),
    .A2(\simon1.seq[19][1] ),
    .A1(net66));
 sg13g2_nor2b_1 _1812_ (.A(net69),
    .B_N(\simon1.seq[1][1] ),
    .Y(_0684_));
 sg13g2_nand2b_2 _1813_ (.Y(_0685_),
    .B(net71),
    .A_N(_0004_));
 sg13g2_a22oi_1 _1814_ (.Y(_0686_),
    .B1(_0684_),
    .B2(_0685_),
    .A2(\simon1.seq[3][1] ),
    .A1(net69));
 sg13g2_nor2b_1 _1815_ (.A(net67),
    .B_N(\simon1.seq[16][1] ),
    .Y(_0687_));
 sg13g2_nand2b_2 _1816_ (.Y(_0688_),
    .B(_0004_),
    .A_N(net71));
 sg13g2_a22oi_1 _1817_ (.Y(_0689_),
    .B1(_0687_),
    .B2(_0688_),
    .A2(\simon1.seq[18][1] ),
    .A1(net67));
 sg13g2_or2_1 _1818_ (.X(_0690_),
    .B(_0004_),
    .A(net71));
 sg13g2_buf_1 fanout84 (.A(net86),
    .X(net84));
 sg13g2_mux2_1 _1820_ (.A0(\simon1.seq[0][1] ),
    .A1(\simon1.seq[2][1] ),
    .S(net70),
    .X(_0692_));
 sg13g2_nor2_1 _1821_ (.A(_0002_),
    .B(_0003_),
    .Y(_0693_));
 sg13g2_o21ai_1 _1822_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_0690_),
    .A2(_0692_));
 sg13g2_or4_1 _1823_ (.A(_0683_),
    .B(_0686_),
    .C(_0689_),
    .D(_0694_),
    .X(_0695_));
 sg13g2_nor2b_1 _1824_ (.A(net69),
    .B_N(\simon1.seq[21][1] ),
    .Y(_0696_));
 sg13g2_a22oi_1 _1825_ (.Y(_0697_),
    .B1(_0681_),
    .B2(_0696_),
    .A2(\simon1.seq[23][1] ),
    .A1(net69));
 sg13g2_nor2b_1 _1826_ (.A(net65),
    .B_N(\simon1.seq[5][1] ),
    .Y(_0698_));
 sg13g2_a22oi_1 _1827_ (.Y(_0699_),
    .B1(_0685_),
    .B2(_0698_),
    .A2(\simon1.seq[7][1] ),
    .A1(net65));
 sg13g2_nor2b_1 _1828_ (.A(net65),
    .B_N(\simon1.seq[20][1] ),
    .Y(_0700_));
 sg13g2_a22oi_1 _1829_ (.Y(_0701_),
    .B1(_0688_),
    .B2(_0700_),
    .A2(\simon1.seq[22][1] ),
    .A1(net65));
 sg13g2_mux2_1 _1830_ (.A0(\simon1.seq[4][1] ),
    .A1(\simon1.seq[6][1] ),
    .S(net67),
    .X(_0702_));
 sg13g2_nor2b_1 _1831_ (.A(_0003_),
    .B_N(_0002_),
    .Y(_0703_));
 sg13g2_o21ai_1 _1832_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0690_),
    .A2(_0702_));
 sg13g2_or4_1 _1833_ (.A(_0697_),
    .B(_0699_),
    .C(_0701_),
    .D(_0704_),
    .X(_0705_));
 sg13g2_nand4_1 _1834_ (.B(_0679_),
    .C(_0695_),
    .A(_0673_),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_buf_2 fanout83 (.A(net86),
    .X(net83));
 sg13g2_xor2_1 _1836_ (.B(_0706_),
    .A(\simon1.user_input[1] ),
    .X(_0708_));
 sg13g2_buf_2 fanout82 (.A(net1),
    .X(net82));
 sg13g2_mux4_1 _1838_ (.S0(net71),
    .A0(\simon1.seq[12][0] ),
    .A1(\simon1.seq[13][0] ),
    .A2(\simon1.seq[14][0] ),
    .A3(\simon1.seq[15][0] ),
    .S1(net68),
    .X(_0710_));
 sg13g2_mux4_1 _1839_ (.S0(net72),
    .A0(\simon1.seq[28][0] ),
    .A1(\simon1.seq[29][0] ),
    .A2(\simon1.seq[30][0] ),
    .A3(\simon1.seq[31][0] ),
    .S1(net70),
    .X(_0711_));
 sg13g2_mux2_1 _1840_ (.A0(_0710_),
    .A1(_0711_),
    .S(_0004_),
    .X(_0712_));
 sg13g2_nand3_1 _1841_ (.B(_0003_),
    .C(_0712_),
    .A(_0002_),
    .Y(_0713_));
 sg13g2_mux4_1 _1842_ (.S0(net71),
    .A0(\simon1.seq[8][0] ),
    .A1(\simon1.seq[9][0] ),
    .A2(\simon1.seq[10][0] ),
    .A3(\simon1.seq[11][0] ),
    .S1(net68),
    .X(_0714_));
 sg13g2_mux4_1 _1843_ (.S0(net72),
    .A0(\simon1.seq[24][0] ),
    .A1(\simon1.seq[25][0] ),
    .A2(\simon1.seq[26][0] ),
    .A3(\simon1.seq[27][0] ),
    .S1(net70),
    .X(_0715_));
 sg13g2_mux2_1 _1844_ (.A0(_0714_),
    .A1(_0715_),
    .S(_0004_),
    .X(_0716_));
 sg13g2_nand2_1 _1845_ (.Y(_0717_),
    .A(_0674_),
    .B(_0716_));
 sg13g2_nor2b_1 _1846_ (.A(net66),
    .B_N(\simon1.seq[17][0] ),
    .Y(_0718_));
 sg13g2_a22oi_1 _1847_ (.Y(_0719_),
    .B1(_0681_),
    .B2(_0718_),
    .A2(\simon1.seq[19][0] ),
    .A1(net66));
 sg13g2_nor2b_1 _1848_ (.A(net69),
    .B_N(\simon1.seq[1][0] ),
    .Y(_0720_));
 sg13g2_a22oi_1 _1849_ (.Y(_0721_),
    .B1(_0685_),
    .B2(_0720_),
    .A2(net69),
    .A1(\simon1.seq[3][0] ));
 sg13g2_nor2b_1 _1850_ (.A(net67),
    .B_N(\simon1.seq[16][0] ),
    .Y(_0722_));
 sg13g2_a22oi_1 _1851_ (.Y(_0723_),
    .B1(_0688_),
    .B2(_0722_),
    .A2(\simon1.seq[18][0] ),
    .A1(net67));
 sg13g2_mux2_1 _1852_ (.A0(\simon1.seq[0][0] ),
    .A1(\simon1.seq[2][0] ),
    .S(net70),
    .X(_0724_));
 sg13g2_o21ai_1 _1853_ (.B1(_0693_),
    .Y(_0725_),
    .A1(_0690_),
    .A2(_0724_));
 sg13g2_or4_1 _1854_ (.A(_0719_),
    .B(_0721_),
    .C(_0723_),
    .D(_0725_),
    .X(_0726_));
 sg13g2_nor2b_1 _1855_ (.A(net69),
    .B_N(\simon1.seq[21][0] ),
    .Y(_0727_));
 sg13g2_a22oi_1 _1856_ (.Y(_0728_),
    .B1(_0681_),
    .B2(_0727_),
    .A2(\simon1.seq[23][0] ),
    .A1(net69));
 sg13g2_nor2b_1 _1857_ (.A(net65),
    .B_N(\simon1.seq[5][0] ),
    .Y(_0729_));
 sg13g2_a22oi_1 _1858_ (.Y(_0730_),
    .B1(_0685_),
    .B2(_0729_),
    .A2(\simon1.seq[7][0] ),
    .A1(net65));
 sg13g2_nor2b_1 _1859_ (.A(net65),
    .B_N(\simon1.seq[20][0] ),
    .Y(_0731_));
 sg13g2_a22oi_1 _1860_ (.Y(_0732_),
    .B1(_0688_),
    .B2(_0731_),
    .A2(\simon1.seq[22][0] ),
    .A1(net65));
 sg13g2_mux2_1 _1861_ (.A0(\simon1.seq[4][0] ),
    .A1(\simon1.seq[6][0] ),
    .S(net67),
    .X(_0733_));
 sg13g2_o21ai_1 _1862_ (.B1(_0703_),
    .Y(_0734_),
    .A1(_0690_),
    .A2(_0733_));
 sg13g2_or4_1 _1863_ (.A(_0728_),
    .B(_0730_),
    .C(_0732_),
    .D(_0734_),
    .X(_0735_));
 sg13g2_nand4_1 _1864_ (.B(_0717_),
    .C(_0726_),
    .A(_0713_),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_buf_2 fanout81 (.A(net82),
    .X(net81));
 sg13g2_xor2_1 _1866_ (.B(net41),
    .A(\simon1.user_input[0] ),
    .X(_0738_));
 sg13g2_nor2_1 _1867_ (.A(_0708_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_buf_2 fanout80 (.A(net82),
    .X(net80));
 sg13g2_buf_1 fanout79 (.A(_0754_),
    .X(net79));
 sg13g2_nor2_1 _1870_ (.A(\simon1.millis_counter[1] ),
    .B(net64),
    .Y(_0742_));
 sg13g2_inv_1 _1871_ (.Y(_0743_),
    .A(\simon1.millis_counter[8] ));
 sg13g2_nor2_1 _1872_ (.A(\simon1.millis_counter[9] ),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand3_1 _1873_ (.B(_0742_),
    .C(_0744_),
    .A(\simon1.millis_counter[2] ),
    .Y(_0745_));
 sg13g2_buf_2 fanout78 (.A(net79),
    .X(net78));
 sg13g2_buf_2 fanout77 (.A(net78),
    .X(net77));
 sg13g2_nand3b_1 _1876_ (.B(\simon1.millis_counter[5] ),
    .C(\simon1.millis_counter[3] ),
    .Y(_0748_),
    .A_N(\simon1.millis_counter[4] ));
 sg13g2_nor4_1 _1877_ (.A(\simon1.millis_counter[7] ),
    .B(\simon1.millis_counter[6] ),
    .C(_0745_),
    .D(_0748_),
    .Y(_0749_));
 sg13g2_buf_2 fanout76 (.A(net79),
    .X(net76));
 sg13g2_buf_2 fanout75 (.A(_0754_),
    .X(net75));
 sg13g2_buf_2 fanout74 (.A(net75),
    .X(net74));
 sg13g2_nand3b_1 _1881_ (.B(net40),
    .C(net57),
    .Y(_0753_),
    .A_N(_0739_));
 sg13g2_inv_1 _1882_ (.Y(_0754_),
    .A(net80));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout72 (.A(_0000_),
    .X(net72));
 sg13g2_a21oi_1 _1885_ (.A1(_0663_),
    .A2(_0753_),
    .Y(_0012_),
    .B1(net76));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(_0000_));
 sg13g2_inv_1 _1887_ (.Y(_0758_),
    .A(\simon1.millis_counter[7] ));
 sg13g2_nand2b_1 _1888_ (.Y(_0759_),
    .B(\simon1.millis_counter[4] ),
    .A_N(\simon1.millis_counter[5] ));
 sg13g2_nor4_2 _1889_ (.A(\simon1.millis_counter[3] ),
    .B(_0758_),
    .C(\simon1.millis_counter[6] ),
    .Y(_0760_),
    .D(_0759_));
 sg13g2_nor3_1 _1890_ (.A(\simon1.millis_counter[1] ),
    .B(net64),
    .C(\simon1.millis_counter[2] ),
    .Y(_0761_));
 sg13g2_nand3_1 _1891_ (.B(_0760_),
    .C(_0761_),
    .A(_0744_),
    .Y(_0762_));
 sg13g2_and2_1 _1892_ (.A(net54),
    .B(_0762_),
    .X(_0763_));
 sg13g2_o21ai_1 _1893_ (.B1(net84),
    .Y(_0764_),
    .A1(\simon1.state[2] ),
    .A2(_0763_));
 sg13g2_inv_1 _1894_ (.Y(_0011_),
    .A(_0764_));
 sg13g2_xor2_1 _1895_ (.B(net5),
    .A(net4),
    .X(_0765_));
 sg13g2_o21ai_1 _1896_ (.B1(net3),
    .Y(_0766_),
    .A1(net4),
    .A2(net5));
 sg13g2_o21ai_1 _1897_ (.B1(_0766_),
    .Y(_0767_),
    .A1(net3),
    .A2(_0765_));
 sg13g2_nand3b_1 _1898_ (.B(_0655_),
    .C(net2),
    .Y(_0768_),
    .A_N(net3));
 sg13g2_o21ai_1 _1899_ (.B1(_0768_),
    .Y(_0769_),
    .A1(net2),
    .A2(_0767_));
 sg13g2_nand3_1 _1900_ (.B(\simon1.state[1] ),
    .C(_0769_),
    .A(net85),
    .Y(_0770_));
 sg13g2_inv_1 _1901_ (.Y(_0771_),
    .A(net55));
 sg13g2_nor2_2 _1902_ (.A(_0771_),
    .B(net40),
    .Y(_0772_));
 sg13g2_nand2_1 _1903_ (.Y(_0773_),
    .A(net86),
    .B(_0772_));
 sg13g2_nand2_1 _1904_ (.Y(_0010_),
    .A(_0770_),
    .B(_0773_));
 sg13g2_nand2_1 _1905_ (.Y(_0774_),
    .A(\simon1.millis_counter[7] ),
    .B(\simon1.millis_counter[6] ));
 sg13g2_nand2_1 _1906_ (.Y(_0775_),
    .A(\simon1.millis_counter[4] ),
    .B(\simon1.millis_counter[5] ));
 sg13g2_nor4_1 _1907_ (.A(\simon1.millis_counter[3] ),
    .B(_0745_),
    .C(_0774_),
    .D(_0775_),
    .Y(_0776_));
 sg13g2_nand2b_1 _1908_ (.Y(_0777_),
    .B(\simon1.state[4] ),
    .A_N(_0776_));
 sg13g2_o21ai_1 _1909_ (.B1(_0657_),
    .Y(_0778_),
    .A1(\simon1.state[0] ),
    .A2(\simon1.state[7] ));
 sg13g2_a21oi_1 _1910_ (.A1(_0777_),
    .A2(_0778_),
    .Y(_0009_),
    .B1(net76));
 sg13g2_buf_2 fanout70 (.A(_0001_),
    .X(net70));
 sg13g2_nor2_1 _1912_ (.A(\simon1.millis_counter[9] ),
    .B(\simon1.millis_counter[8] ),
    .Y(_0780_));
 sg13g2_nor2b_1 _1913_ (.A(net64),
    .B_N(\simon1.millis_counter[1] ),
    .Y(_0781_));
 sg13g2_nand4_1 _1914_ (.B(_0760_),
    .C(_0780_),
    .A(\simon1.millis_counter[2] ),
    .Y(_0782_),
    .D(_0781_));
 sg13g2_buf_2 fanout69 (.A(net70),
    .X(net69));
 sg13g2_nand2_1 _1916_ (.Y(_0784_),
    .A(net52),
    .B(net50));
 sg13g2_nor3_1 _1917_ (.A(net47),
    .B(_0782_),
    .C(_0784_),
    .Y(_0785_));
 sg13g2_buf_2 fanout68 (.A(_0001_),
    .X(net68));
 sg13g2_nand2b_1 _1919_ (.Y(_0787_),
    .B(net58),
    .A_N(_0785_));
 sg13g2_inv_1 _1920_ (.Y(_0788_),
    .A(_0029_));
 sg13g2_buf_2 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_1 fanout66 (.A(net67),
    .X(net66));
 sg13g2_nand2_2 _1923_ (.Y(_0791_),
    .A(\simon1.seq_counter[0] ),
    .B(\simon1.seq_counter[1] ));
 sg13g2_a22oi_1 _1924_ (.Y(_0792_),
    .B1(_0791_),
    .B2(_0788_),
    .A2(\simon1.seq_counter[4] ),
    .A1(\simon1.seq_counter[3] ));
 sg13g2_a21oi_1 _1925_ (.A1(_0788_),
    .A2(_0791_),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_inv_1 _1926_ (.Y(_0794_),
    .A(\simon1.seq_counter[3] ));
 sg13g2_and3_1 _1927_ (.X(_0795_),
    .A(\simon1.seq_counter[0] ),
    .B(\simon1.seq_counter[1] ),
    .C(\simon1.seq_counter[2] ));
 sg13g2_buf_2 fanout65 (.A(net67),
    .X(net65));
 sg13g2_nor3_1 _1929_ (.A(_0794_),
    .B(_0030_),
    .C(_0795_),
    .Y(_0797_));
 sg13g2_xnor2_1 _1930_ (.Y(_0798_),
    .A(_0030_),
    .B(_0795_));
 sg13g2_nor2_1 _1931_ (.A(\simon1.seq_counter[3] ),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_xor2_1 _1932_ (.B(_0031_),
    .A(\simon1.seq_counter[4] ),
    .X(_0800_));
 sg13g2_o21ai_1 _1933_ (.B1(_0800_),
    .Y(_0801_),
    .A1(_0797_),
    .A2(_0799_));
 sg13g2_and2_1 _1934_ (.A(\simon1.seq_counter[3] ),
    .B(_0795_),
    .X(_0802_));
 sg13g2_nand3b_1 _1935_ (.B(_0802_),
    .C(_0030_),
    .Y(_0803_),
    .A_N(_0031_));
 sg13g2_xnor2_1 _1936_ (.Y(_0804_),
    .A(_0029_),
    .B(_0791_));
 sg13g2_xor2_1 _1937_ (.B(_0028_),
    .A(\simon1.seq_counter[1] ),
    .X(_0805_));
 sg13g2_buf_2 fanout64 (.A(\simon1.millis_counter[0] ),
    .X(net64));
 sg13g2_nand2b_1 _1939_ (.Y(_0807_),
    .B(\simon1.seq_counter[0] ),
    .A_N(net60));
 sg13g2_inv_1 _1940_ (.Y(_0808_),
    .A(\simon1.seq_counter[0] ));
 sg13g2_nand3_1 _1941_ (.B(_0808_),
    .C(_0805_),
    .A(net59),
    .Y(_0809_));
 sg13g2_o21ai_1 _1942_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0805_),
    .A2(_0807_));
 sg13g2_o21ai_1 _1943_ (.B1(_0810_),
    .Y(_0811_),
    .A1(\simon1.seq_counter[2] ),
    .A2(_0804_));
 sg13g2_a221oi_1 _1944_ (.B2(_0803_),
    .C1(_0811_),
    .B1(_0801_),
    .A1(\simon1.seq_counter[2] ),
    .Y(_0812_),
    .A2(_0793_));
 sg13g2_buf_2 fanout63 (.A(\simon1.play1.freq[3] ),
    .X(net63));
 sg13g2_or4_2 _1946_ (.A(\simon1.millis_counter[7] ),
    .B(\simon1.millis_counter[6] ),
    .C(_0745_),
    .D(_0748_),
    .X(_0814_));
 sg13g2_buf_2 fanout62 (.A(\simon1.play1.freq[6] ),
    .X(net62));
 sg13g2_nor3_1 _1948_ (.A(_0708_),
    .B(_0738_),
    .C(_0814_),
    .Y(_0816_));
 sg13g2_buf_2 fanout61 (.A(\simon1.score1.active_digit ),
    .X(net61));
 sg13g2_nand3_1 _1950_ (.B(net39),
    .C(_0816_),
    .A(net56),
    .Y(_0818_));
 sg13g2_a21oi_1 _1951_ (.A1(_0787_),
    .A2(_0818_),
    .Y(_0008_),
    .B1(net76));
 sg13g2_nand4_1 _1952_ (.B(_0744_),
    .C(_0760_),
    .A(net54),
    .Y(_0819_),
    .D(_0761_));
 sg13g2_nand2_1 _1953_ (.Y(_0820_),
    .A(net58),
    .B(_0785_));
 sg13g2_o21ai_1 _1954_ (.B1(_0820_),
    .Y(_0821_),
    .A1(net39),
    .A2(_0819_));
 sg13g2_buf_1 fanout60 (.A(\simon1.seq_length[0] ),
    .X(net60));
 sg13g2_and3_1 _1956_ (.X(_0089_),
    .A(\simon1.state[4] ),
    .B(net84),
    .C(_0776_));
 sg13g2_a21o_1 _1957_ (.A2(_0821_),
    .A1(net84),
    .B1(_0089_),
    .X(_0007_));
 sg13g2_inv_1 _1958_ (.Y(_0823_),
    .A(\simon1.state[1] ));
 sg13g2_nand2_1 _1959_ (.Y(_0824_),
    .A(net56),
    .B(_0816_));
 sg13g2_mux2_1 _1960_ (.A0(_0824_),
    .A1(_0819_),
    .S(net39),
    .X(_0825_));
 sg13g2_o21ai_1 _1961_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_0823_),
    .A2(_0769_));
 sg13g2_and2_1 _1962_ (.A(net86),
    .B(_0826_),
    .X(_0006_));
 sg13g2_buf_2 fanout59 (.A(\simon1.seq_length[0] ),
    .X(net59));
 sg13g2_buf_2 fanout58 (.A(\simon1.state[3] ),
    .X(net58));
 sg13g2_xor2_1 _1965_ (.B(net6),
    .A(\simon1.score1.active_digit ),
    .X(_0015_));
 sg13g2_inv_1 _1966_ (.Y(_0014_),
    .A(_0015_));
 sg13g2_buf_2 fanout57 (.A(\simon1.state[5] ),
    .X(net57));
 sg13g2_inv_1 _1968_ (.Y(_0830_),
    .A(\simon1.score1.ena ));
 sg13g2_buf_1 fanout56 (.A(net57),
    .X(net56));
 sg13g2_nor2b_1 _1970_ (.A(net61),
    .B_N(\simon1.score1.ones[1] ),
    .Y(_0832_));
 sg13g2_a22oi_1 _1971_ (.Y(_0833_),
    .B1(_0830_),
    .B2(_0832_),
    .A2(\simon1.score1.tens[1] ),
    .A1(net61));
 sg13g2_inv_1 _1972_ (.Y(_0834_),
    .A(_0833_));
 sg13g2_inv_1 _1973_ (.Y(_0835_),
    .A(\simon1.score1.ones[2] ));
 sg13g2_nor2_1 _1974_ (.A(_0835_),
    .B(net61),
    .Y(_0836_));
 sg13g2_a22oi_1 _1975_ (.Y(_0837_),
    .B1(_0027_),
    .B2(_0836_),
    .A2(\simon1.score1.tens[2] ),
    .A1(net61));
 sg13g2_buf_2 fanout55 (.A(net57),
    .X(net55));
 sg13g2_nand2b_1 _1977_ (.Y(_0839_),
    .B(\simon1.score1.ones[0] ),
    .A_N(net61));
 sg13g2_nand2_1 _1978_ (.Y(_0840_),
    .A(net61),
    .B(\simon1.score1.tens[0] ));
 sg13g2_nand3_1 _1979_ (.B(_0839_),
    .C(_0840_),
    .A(\simon1.score1.ena ),
    .Y(_0841_));
 sg13g2_buf_2 fanout54 (.A(\simon1.state[6] ),
    .X(net54));
 sg13g2_nor2_1 _1981_ (.A(_0837_),
    .B(_0841_),
    .Y(_0843_));
 sg13g2_inv_1 _1982_ (.Y(_0844_),
    .A(\simon1.score1.ones[3] ));
 sg13g2_nor2_1 _1983_ (.A(_0844_),
    .B(net61),
    .Y(_0845_));
 sg13g2_a22oi_1 _1984_ (.Y(_0846_),
    .B1(_0027_),
    .B2(_0845_),
    .A2(\simon1.score1.tens[3] ),
    .A1(net61));
 sg13g2_buf_1 fanout53 (.A(\simon1.tone_sequence_counter[0] ),
    .X(net53));
 sg13g2_nand3_1 _1986_ (.B(_0837_),
    .C(_0841_),
    .A(_0846_),
    .Y(_0848_));
 sg13g2_nor2b_1 _1987_ (.A(_0843_),
    .B_N(_0848_),
    .Y(_0849_));
 sg13g2_inv_1 _1988_ (.Y(_0850_),
    .A(_0837_));
 sg13g2_nor2_1 _1989_ (.A(_0834_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_or2_1 _1990_ (.X(_0852_),
    .B(_0851_),
    .A(_0846_));
 sg13g2_buf_2 fanout52 (.A(\simon1.tone_sequence_counter[0] ),
    .X(net52));
 sg13g2_o21ai_1 _1992_ (.B1(_0852_),
    .Y(_0854_),
    .A1(_0834_),
    .A2(_0849_));
 sg13g2_xnor2_1 _1993_ (.Y(_0204_),
    .A(net6),
    .B(_0854_));
 sg13g2_xor2_1 _1994_ (.B(_0841_),
    .A(_0833_),
    .X(_0855_));
 sg13g2_o21ai_1 _1995_ (.B1(_0852_),
    .Y(_0856_),
    .A1(_0837_),
    .A2(_0855_));
 sg13g2_xnor2_1 _1996_ (.Y(_0205_),
    .A(net6),
    .B(_0856_));
 sg13g2_o21ai_1 _1997_ (.B1(_0846_),
    .Y(_0857_),
    .A1(_0850_),
    .A2(_0841_));
 sg13g2_nor2b_1 _1998_ (.A(_0851_),
    .B_N(_0857_),
    .Y(_0858_));
 sg13g2_xnor2_1 _1999_ (.Y(_0206_),
    .A(net6),
    .B(_0858_));
 sg13g2_nor2_1 _2000_ (.A(_0833_),
    .B(_0837_),
    .Y(_0859_));
 sg13g2_nand2_1 _2001_ (.Y(_0860_),
    .A(_0846_),
    .B(_0851_));
 sg13g2_nand2b_1 _2002_ (.Y(_0861_),
    .B(_0860_),
    .A_N(_0859_));
 sg13g2_inv_1 _2003_ (.Y(_0862_),
    .A(_0852_));
 sg13g2_a221oi_1 _2004_ (.B2(_0841_),
    .C1(_0862_),
    .B1(_0861_),
    .A1(_0833_),
    .Y(_0863_),
    .A2(_0843_));
 sg13g2_xor2_1 _2005_ (.B(_0863_),
    .A(net6),
    .X(_0207_));
 sg13g2_a21oi_1 _2006_ (.A1(_0846_),
    .A2(_0834_),
    .Y(_0864_),
    .B1(_0851_));
 sg13g2_nor2_1 _2007_ (.A(_0841_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_xor2_1 _2008_ (.B(_0865_),
    .A(net6),
    .X(_0208_));
 sg13g2_a21o_1 _2009_ (.A2(_0837_),
    .A1(_0846_),
    .B1(_0834_),
    .X(_0866_));
 sg13g2_a21oi_1 _2010_ (.A1(_0846_),
    .A2(_0850_),
    .Y(_0867_),
    .B1(_0851_));
 sg13g2_a21oi_1 _2011_ (.A1(_0841_),
    .A2(_0866_),
    .Y(_0868_),
    .B1(_0867_));
 sg13g2_xor2_1 _2012_ (.B(_0868_),
    .A(net6),
    .X(_0209_));
 sg13g2_nand2_1 _2013_ (.Y(_0869_),
    .A(_0841_),
    .B(_0859_));
 sg13g2_nand3_1 _2014_ (.B(_0860_),
    .C(_0869_),
    .A(_0852_),
    .Y(_0870_));
 sg13g2_xnor2_1 _2015_ (.Y(_0210_),
    .A(net6),
    .B(_0870_));
 sg13g2_buf_2 fanout51 (.A(\simon1.tone_sequence_counter[1] ),
    .X(net51));
 sg13g2_inv_1 _2017_ (.Y(_0872_),
    .A(_0035_));
 sg13g2_inv_2 _2018_ (.Y(_0873_),
    .A(net58));
 sg13g2_nor2_1 _2019_ (.A(\simon1.state[4] ),
    .B(net56),
    .Y(_0874_));
 sg13g2_nand3b_1 _2020_ (.B(_0873_),
    .C(_0874_),
    .Y(_0875_),
    .A_N(net54));
 sg13g2_or2_1 _2021_ (.X(_0876_),
    .B(_0875_),
    .A(\simon1.state[2] ));
 sg13g2_a21oi_1 _2022_ (.A1(\simon1.state[0] ),
    .A2(\simon1.state[1] ),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_o21ai_1 _2023_ (.B1(_0657_),
    .Y(_0878_),
    .A1(_0872_),
    .A2(_0877_));
 sg13g2_inv_1 _2024_ (.Y(_0879_),
    .A(_0028_));
 sg13g2_nand4_1 _2025_ (.B(_0654_),
    .C(_0035_),
    .A(net84),
    .Y(_0880_),
    .D(_0657_));
 sg13g2_nor2_2 _2026_ (.A(_0876_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_o21ai_1 _2027_ (.B1(_0881_),
    .Y(_0882_),
    .A1(net59),
    .A2(_0879_));
 sg13g2_buf_2 fanout50 (.A(\simon1.tone_sequence_counter[1] ),
    .X(net50));
 sg13g2_or2_1 _2029_ (.X(_0884_),
    .B(\simon1.seq_length[2] ),
    .A(\simon1.seq_length[3] ));
 sg13g2_o21ai_1 _2030_ (.B1(_0881_),
    .Y(_0885_),
    .A1(\simon1.seq_length[4] ),
    .A2(_0884_));
 sg13g2_nand2_1 _2031_ (.Y(_0886_),
    .A(_0882_),
    .B(_0885_));
 sg13g2_nor2_1 _2032_ (.A(_0878_),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_and2_1 _2033_ (.A(\simon1.seq[0][0] ),
    .B(_0878_),
    .X(_0888_));
 sg13g2_a21oi_1 _2034_ (.A1(\simon1.next_random[0] ),
    .A2(_0887_),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_nand2_1 _2035_ (.Y(_0890_),
    .A(\simon1.seq[0][0] ),
    .B(_0886_));
 sg13g2_o21ai_1 _2036_ (.B1(_0890_),
    .Y(_0038_),
    .A1(net75),
    .A2(_0889_));
 sg13g2_inv_1 _2037_ (.Y(_0891_),
    .A(_0878_));
 sg13g2_and3_1 _2038_ (.X(_0892_),
    .A(net81),
    .B(\simon1.next_random[1] ),
    .C(_0891_));
 sg13g2_buf_2 fanout49 (.A(\simon1.tone_sequence_counter[2] ),
    .X(net49));
 sg13g2_buf_2 fanout48 (.A(net49),
    .X(net48));
 sg13g2_nand2b_2 _2041_ (.Y(_0895_),
    .B(_0881_),
    .A_N(\simon1.seq_length[4] ));
 sg13g2_nand2b_1 _2042_ (.Y(_0896_),
    .B(\simon1.seq_length[3] ),
    .A_N(\simon1.seq_length[2] ));
 sg13g2_nor2_1 _2043_ (.A(_0895_),
    .B(_0896_),
    .Y(_0897_));
 sg13g2_and2_1 _2044_ (.A(_0882_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_mux2_1 _2045_ (.A0(\simon1.seq[8][1] ),
    .A1(net28),
    .S(_0898_),
    .X(_0039_));
 sg13g2_buf_2 fanout47 (.A(_0033_),
    .X(net47));
 sg13g2_nand2_1 _2047_ (.Y(_0900_),
    .A(\simon1.seq_length[3] ),
    .B(\simon1.seq_length[2] ));
 sg13g2_or2_1 _2048_ (.X(_0901_),
    .B(_0900_),
    .A(_0895_));
 sg13g2_buf_2 fanout46 (.A(_0998_),
    .X(net46));
 sg13g2_buf_2 fanout45 (.A(_1075_),
    .X(net45));
 sg13g2_and2_1 _2051_ (.A(_0879_),
    .B(_0881_),
    .X(_0904_));
 sg13g2_nor2b_2 _2052_ (.A(net59),
    .B_N(_0904_),
    .Y(_0905_));
 sg13g2_nand2b_1 _2053_ (.Y(_0906_),
    .B(_0905_),
    .A_N(_0901_));
 sg13g2_mux2_1 _2054_ (.A0(net28),
    .A1(\simon1.seq[14][1] ),
    .S(_0906_),
    .X(_0040_));
 sg13g2_nand3_1 _2055_ (.B(_0028_),
    .C(_0881_),
    .A(net59),
    .Y(_0907_));
 sg13g2_nor2_1 _2056_ (.A(_0901_),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_mux2_1 _2057_ (.A0(\simon1.seq[13][1] ),
    .A1(net28),
    .S(_0908_),
    .X(_0041_));
 sg13g2_nor2b_1 _2058_ (.A(_0901_),
    .B_N(_0882_),
    .Y(_0909_));
 sg13g2_mux2_1 _2059_ (.A0(\simon1.seq[12][1] ),
    .A1(net28),
    .S(_0909_),
    .X(_0042_));
 sg13g2_and3_1 _2060_ (.X(_0910_),
    .A(net81),
    .B(\simon1.next_random[0] ),
    .C(_0891_));
 sg13g2_buf_2 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_1 fanout43 (.A(_0227_),
    .X(net43));
 sg13g2_and2_1 _2063_ (.A(net59),
    .B(_0904_),
    .X(_0913_));
 sg13g2_buf_2 fanout42 (.A(_0227_),
    .X(net42));
 sg13g2_nand2_1 _2065_ (.Y(_0915_),
    .A(_0885_),
    .B(_0913_));
 sg13g2_mux2_1 _2066_ (.A0(net27),
    .A1(\simon1.seq[3][0] ),
    .S(_0915_),
    .X(_0043_));
 sg13g2_buf_2 fanout41 (.A(_0736_),
    .X(net41));
 sg13g2_nand2_1 _2068_ (.Y(_0917_),
    .A(net59),
    .B(_0904_));
 sg13g2_and2_1 _2069_ (.A(\simon1.seq_length[4] ),
    .B(_0881_),
    .X(_0918_));
 sg13g2_nand2b_1 _2070_ (.Y(_0919_),
    .B(_0918_),
    .A_N(_0900_));
 sg13g2_nor2_1 _2071_ (.A(_0917_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_mux2_1 _2072_ (.A0(\simon1.seq[31][0] ),
    .A1(net26),
    .S(_0920_),
    .X(_0044_));
 sg13g2_and2_1 _2073_ (.A(_0885_),
    .B(_0905_),
    .X(_0921_));
 sg13g2_mux2_1 _2074_ (.A0(\simon1.seq[2][0] ),
    .A1(net27),
    .S(_0921_),
    .X(_0045_));
 sg13g2_and3_1 _2075_ (.X(_0922_),
    .A(net59),
    .B(_0028_),
    .C(_0881_));
 sg13g2_buf_2 fanout40 (.A(_0749_),
    .X(net40));
 sg13g2_nand2_2 _2077_ (.Y(_0924_),
    .A(\simon1.seq_length[4] ),
    .B(_0881_));
 sg13g2_nor2_1 _2078_ (.A(_0900_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nand2_1 _2079_ (.Y(_0926_),
    .A(_0922_),
    .B(_0925_));
 sg13g2_mux2_1 _2080_ (.A0(net26),
    .A1(\simon1.seq[29][0] ),
    .S(_0926_),
    .X(_0046_));
 sg13g2_nand2_1 _2081_ (.Y(_0927_),
    .A(_0882_),
    .B(_0925_));
 sg13g2_mux2_1 _2082_ (.A0(net26),
    .A1(\simon1.seq[28][0] ),
    .S(_0927_),
    .X(_0047_));
 sg13g2_nand2b_1 _2083_ (.Y(_0928_),
    .B(_0918_),
    .A_N(_0896_));
 sg13g2_nor2_1 _2084_ (.A(_0917_),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_mux2_1 _2085_ (.A0(\simon1.seq[27][0] ),
    .A1(net26),
    .S(_0929_),
    .X(_0048_));
 sg13g2_nand2b_1 _2086_ (.Y(_0930_),
    .B(_0904_),
    .A_N(net59));
 sg13g2_nor2_1 _2087_ (.A(_0930_),
    .B(_0928_),
    .Y(_0931_));
 sg13g2_mux2_1 _2088_ (.A0(\simon1.seq[26][0] ),
    .A1(net26),
    .S(_0931_),
    .X(_0049_));
 sg13g2_nor2_1 _2089_ (.A(_0896_),
    .B(_0924_),
    .Y(_0932_));
 sg13g2_nand2_1 _2090_ (.Y(_0933_),
    .A(_0922_),
    .B(_0932_));
 sg13g2_mux2_1 _2091_ (.A0(net23),
    .A1(\simon1.seq[25][0] ),
    .S(_0933_),
    .X(_0050_));
 sg13g2_nand2_1 _2092_ (.Y(_0934_),
    .A(_0882_),
    .B(_0932_));
 sg13g2_mux2_1 _2093_ (.A0(net26),
    .A1(\simon1.seq[24][0] ),
    .S(_0934_),
    .X(_0051_));
 sg13g2_buf_2 fanout39 (.A(_0812_),
    .X(net39));
 sg13g2_nand2b_1 _2095_ (.Y(_0936_),
    .B(\simon1.seq_length[2] ),
    .A_N(\simon1.seq_length[3] ));
 sg13g2_or2_1 _2096_ (.X(_0937_),
    .B(_0936_),
    .A(_0924_));
 sg13g2_nor2_1 _2097_ (.A(_0917_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_mux2_1 _2098_ (.A0(\simon1.seq[23][0] ),
    .A1(net27),
    .S(_0938_),
    .X(_0052_));
 sg13g2_nor2_1 _2099_ (.A(_0930_),
    .B(_0937_),
    .Y(_0939_));
 sg13g2_mux2_1 _2100_ (.A0(\simon1.seq[22][0] ),
    .A1(net27),
    .S(_0939_),
    .X(_0053_));
 sg13g2_nand2_1 _2101_ (.Y(_0940_),
    .A(_0897_),
    .B(_0913_));
 sg13g2_mux2_1 _2102_ (.A0(net28),
    .A1(\simon1.seq[11][1] ),
    .S(_0940_),
    .X(_0054_));
 sg13g2_nor2_1 _2103_ (.A(_0924_),
    .B(_0936_),
    .Y(_0941_));
 sg13g2_nand2_1 _2104_ (.Y(_0942_),
    .A(_0922_),
    .B(_0941_));
 sg13g2_mux2_1 _2105_ (.A0(net27),
    .A1(\simon1.seq[21][0] ),
    .S(_0942_),
    .X(_0055_));
 sg13g2_nand2_1 _2106_ (.Y(_0943_),
    .A(_0885_),
    .B(_0922_));
 sg13g2_mux2_1 _2107_ (.A0(net26),
    .A1(\simon1.seq[1][0] ),
    .S(_0943_),
    .X(_0056_));
 sg13g2_nor2_1 _2108_ (.A(_0884_),
    .B(_0924_),
    .Y(_0944_));
 sg13g2_and2_1 _2109_ (.A(_0913_),
    .B(_0944_),
    .X(_0945_));
 sg13g2_mux2_1 _2110_ (.A0(\simon1.seq[19][0] ),
    .A1(net25),
    .S(_0945_),
    .X(_0057_));
 sg13g2_and2_1 _2111_ (.A(_0905_),
    .B(_0944_),
    .X(_0946_));
 sg13g2_mux2_1 _2112_ (.A0(\simon1.seq[18][0] ),
    .A1(net24),
    .S(_0946_),
    .X(_0058_));
 sg13g2_nand2_1 _2113_ (.Y(_0947_),
    .A(_0922_),
    .B(_0944_));
 sg13g2_mux2_1 _2114_ (.A0(net24),
    .A1(\simon1.seq[17][0] ),
    .S(_0947_),
    .X(_0059_));
 sg13g2_nand2_1 _2115_ (.Y(_0948_),
    .A(_0882_),
    .B(_0944_));
 sg13g2_mux2_1 _2116_ (.A0(net24),
    .A1(\simon1.seq[16][0] ),
    .S(_0948_),
    .X(_0060_));
 sg13g2_nand2b_1 _2117_ (.Y(_0949_),
    .B(_0913_),
    .A_N(_0901_));
 sg13g2_mux2_1 _2118_ (.A0(net23),
    .A1(\simon1.seq[15][0] ),
    .S(_0949_),
    .X(_0061_));
 sg13g2_mux2_1 _2119_ (.A0(net23),
    .A1(\simon1.seq[14][0] ),
    .S(_0906_),
    .X(_0062_));
 sg13g2_mux2_1 _2120_ (.A0(\simon1.seq[13][0] ),
    .A1(net23),
    .S(_0908_),
    .X(_0063_));
 sg13g2_nand2_1 _2121_ (.Y(_0950_),
    .A(_0897_),
    .B(_0905_));
 sg13g2_mux2_1 _2122_ (.A0(net28),
    .A1(\simon1.seq[10][1] ),
    .S(_0950_),
    .X(_0064_));
 sg13g2_mux2_1 _2123_ (.A0(\simon1.seq[12][0] ),
    .A1(net23),
    .S(_0909_),
    .X(_0065_));
 sg13g2_mux2_1 _2124_ (.A0(net23),
    .A1(\simon1.seq[11][0] ),
    .S(_0940_),
    .X(_0066_));
 sg13g2_nor3_1 _2125_ (.A(_0895_),
    .B(_0896_),
    .C(_0907_),
    .Y(_0951_));
 sg13g2_mux2_1 _2126_ (.A0(\simon1.seq[9][1] ),
    .A1(net30),
    .S(_0951_),
    .X(_0067_));
 sg13g2_mux2_1 _2127_ (.A0(\simon1.seq[9][0] ),
    .A1(net25),
    .S(_0951_),
    .X(_0068_));
 sg13g2_nor2_1 _2128_ (.A(_0895_),
    .B(_0936_),
    .Y(_0952_));
 sg13g2_nand2_1 _2129_ (.Y(_0953_),
    .A(_0913_),
    .B(_0952_));
 sg13g2_mux2_1 _2130_ (.A0(net29),
    .A1(\simon1.seq[7][1] ),
    .S(_0953_),
    .X(_0069_));
 sg13g2_nand2_1 _2131_ (.Y(_0954_),
    .A(_0905_),
    .B(_0952_));
 sg13g2_mux2_1 _2132_ (.A0(net29),
    .A1(\simon1.seq[6][1] ),
    .S(_0954_),
    .X(_0070_));
 sg13g2_buf_2 fanout38 (.A(_1060_),
    .X(net38));
 sg13g2_nor3_1 _2134_ (.A(_0895_),
    .B(_0907_),
    .C(_0936_),
    .Y(_0956_));
 sg13g2_mux2_1 _2135_ (.A0(\simon1.seq[5][1] ),
    .A1(net29),
    .S(_0956_),
    .X(_0071_));
 sg13g2_mux2_1 _2136_ (.A0(\simon1.seq[8][0] ),
    .A1(net23),
    .S(_0898_),
    .X(_0072_));
 sg13g2_mux2_1 _2137_ (.A0(net24),
    .A1(\simon1.seq[7][0] ),
    .S(_0953_),
    .X(_0073_));
 sg13g2_mux2_1 _2138_ (.A0(net24),
    .A1(\simon1.seq[6][0] ),
    .S(_0954_),
    .X(_0074_));
 sg13g2_mux2_1 _2139_ (.A0(\simon1.seq[5][0] ),
    .A1(net24),
    .S(_0956_),
    .X(_0075_));
 sg13g2_and2_1 _2140_ (.A(_0882_),
    .B(_0952_),
    .X(_0957_));
 sg13g2_mux2_1 _2141_ (.A0(\simon1.seq[4][1] ),
    .A1(net29),
    .S(_0957_),
    .X(_0076_));
 sg13g2_mux2_1 _2142_ (.A0(\simon1.seq[31][1] ),
    .A1(net31),
    .S(_0920_),
    .X(_0077_));
 sg13g2_mux2_1 _2143_ (.A0(net31),
    .A1(\simon1.seq[3][1] ),
    .S(_0915_),
    .X(_0078_));
 sg13g2_mux2_1 _2144_ (.A0(\simon1.seq[4][0] ),
    .A1(net24),
    .S(_0957_),
    .X(_0079_));
 sg13g2_nor2_1 _2145_ (.A(_0930_),
    .B(_0919_),
    .Y(_0958_));
 sg13g2_mux2_1 _2146_ (.A0(\simon1.seq[30][0] ),
    .A1(net26),
    .S(_0958_),
    .X(_0080_));
 sg13g2_mux2_1 _2147_ (.A0(\simon1.seq[30][1] ),
    .A1(net31),
    .S(_0958_),
    .X(_0087_));
 sg13g2_mux2_1 _2148_ (.A0(\simon1.seq[2][1] ),
    .A1(net32),
    .S(_0921_),
    .X(_0088_));
 sg13g2_mux2_1 _2149_ (.A0(net31),
    .A1(\simon1.seq[28][1] ),
    .S(_0927_),
    .X(_0131_));
 sg13g2_xnor2_1 _2150_ (.Y(_0959_),
    .A(net3),
    .B(net5));
 sg13g2_nor4_1 _2151_ (.A(net2),
    .B(net4),
    .C(_0770_),
    .D(_0959_),
    .Y(_0960_));
 sg13g2_a21o_1 _2152_ (.A2(_0770_),
    .A1(\simon1.user_input[0] ),
    .B1(_0960_),
    .X(_0134_));
 sg13g2_and2_1 _2153_ (.A(_0656_),
    .B(_0765_),
    .X(_0961_));
 sg13g2_mux2_1 _2154_ (.A0(_0961_),
    .A1(\simon1.user_input[1] ),
    .S(_0770_),
    .X(_0135_));
 sg13g2_buf_2 fanout37 (.A(_1087_),
    .X(net37));
 sg13g2_inv_1 _2156_ (.Y(_0963_),
    .A(\simon1.state[7] ));
 sg13g2_a21oi_1 _2157_ (.A1(_0873_),
    .A2(_0963_),
    .Y(_0964_),
    .B1(net52));
 sg13g2_buf_2 fanout36 (.A(_1087_),
    .X(net36));
 sg13g2_nor2_2 _2159_ (.A(net52),
    .B(net51),
    .Y(_0966_));
 sg13g2_nand2b_1 _2160_ (.Y(_0967_),
    .B(_0742_),
    .A_N(\simon1.millis_counter[2] ));
 sg13g2_nand2_1 _2161_ (.Y(_0968_),
    .A(\simon1.millis_counter[9] ),
    .B(\simon1.millis_counter[8] ));
 sg13g2_or4_1 _2162_ (.A(_0748_),
    .B(_0967_),
    .C(_0774_),
    .D(_0968_),
    .X(_0969_));
 sg13g2_and3_1 _2163_ (.X(_0970_),
    .A(net48),
    .B(_0966_),
    .C(_0969_));
 sg13g2_nor3_1 _2164_ (.A(net47),
    .B(_0814_),
    .C(_0966_),
    .Y(_0971_));
 sg13g2_o21ai_1 _2165_ (.B1(\simon1.state[7] ),
    .Y(_0972_),
    .A1(_0970_),
    .A2(_0971_));
 sg13g2_nor3_1 _2166_ (.A(\simon1.state[4] ),
    .B(net58),
    .C(_0872_),
    .Y(_0973_));
 sg13g2_and2_1 _2167_ (.A(\simon1.tone_sequence_counter[2] ),
    .B(_0966_),
    .X(_0974_));
 sg13g2_nor3_1 _2168_ (.A(_0035_),
    .B(net40),
    .C(_0974_),
    .Y(_0975_));
 sg13g2_nor2_1 _2169_ (.A(_0973_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_nand2_1 _2170_ (.Y(_0977_),
    .A(net58),
    .B(_0782_));
 sg13g2_and4_1 _2171_ (.A(net85),
    .B(_0972_),
    .C(_0976_),
    .D(_0977_),
    .X(_0978_));
 sg13g2_buf_2 fanout35 (.A(_0816_),
    .X(net35));
 sg13g2_mux2_1 _2173_ (.A0(net52),
    .A1(_0964_),
    .S(_0978_),
    .X(_0138_));
 sg13g2_buf_2 fanout34 (.A(_1063_),
    .X(net34));
 sg13g2_a21oi_1 _2175_ (.A1(_0872_),
    .A2(\simon1.state[7] ),
    .Y(_0981_),
    .B1(net58));
 sg13g2_a21o_1 _2176_ (.A2(net50),
    .A1(net52),
    .B1(_0981_),
    .X(_0982_));
 sg13g2_inv_1 _2177_ (.Y(_0983_),
    .A(net52));
 sg13g2_nand2_1 _2178_ (.Y(_0984_),
    .A(_0872_),
    .B(net49));
 sg13g2_nand2_1 _2179_ (.Y(_0985_),
    .A(_0983_),
    .B(_0984_));
 sg13g2_a21oi_1 _2180_ (.A1(_0978_),
    .A2(_0985_),
    .Y(_0986_),
    .B1(net50));
 sg13g2_a21oi_1 _2181_ (.A1(_0978_),
    .A2(_0982_),
    .Y(_0139_),
    .B1(_0986_));
 sg13g2_buf_2 fanout33 (.A(_0512_),
    .X(net33));
 sg13g2_o21ai_1 _2183_ (.B1(net47),
    .Y(_0988_),
    .A1(net50),
    .A2(_0984_));
 sg13g2_nand3_1 _2184_ (.B(net50),
    .C(net47),
    .A(net52),
    .Y(_0989_));
 sg13g2_o21ai_1 _2185_ (.B1(_0989_),
    .Y(_0990_),
    .A1(net50),
    .A2(net47));
 sg13g2_a21oi_1 _2186_ (.A1(_0983_),
    .A2(_0988_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_nor2_1 _2187_ (.A(_0981_),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_mux2_1 _2188_ (.A0(net49),
    .A1(_0992_),
    .S(_0978_),
    .X(_0140_));
 sg13g2_mux2_1 _2189_ (.A0(\simon1.seq[27][1] ),
    .A1(net30),
    .S(_0929_),
    .X(_0186_));
 sg13g2_mux2_1 _2190_ (.A0(\simon1.seq[18][1] ),
    .A1(net29),
    .S(_0946_),
    .X(_0187_));
 sg13g2_mux2_1 _2191_ (.A0(\simon1.seq[26][1] ),
    .A1(net31),
    .S(_0931_),
    .X(_0188_));
 sg13g2_mux2_1 _2192_ (.A0(net28),
    .A1(\simon1.seq[25][1] ),
    .S(_0933_),
    .X(_0189_));
 sg13g2_mux2_1 _2193_ (.A0(\simon1.seq[22][1] ),
    .A1(net32),
    .S(_0939_),
    .X(_0190_));
 sg13g2_mux2_1 _2194_ (.A0(\simon1.seq[23][1] ),
    .A1(net32),
    .S(_0938_),
    .X(_0191_));
 sg13g2_nand2_1 _2195_ (.Y(_0993_),
    .A(_0882_),
    .B(_0941_));
 sg13g2_mux2_1 _2196_ (.A0(net29),
    .A1(\simon1.seq[20][1] ),
    .S(_0993_),
    .X(_0192_));
 sg13g2_mux2_1 _2197_ (.A0(net31),
    .A1(\simon1.seq[21][1] ),
    .S(_0942_),
    .X(_0193_));
 sg13g2_mux2_1 _2198_ (.A0(net30),
    .A1(\simon1.seq[24][1] ),
    .S(_0934_),
    .X(_0194_));
 sg13g2_mux2_1 _2199_ (.A0(\simon1.seq[19][1] ),
    .A1(net30),
    .S(_0945_),
    .X(_0195_));
 sg13g2_mux2_1 _2200_ (.A0(net29),
    .A1(\simon1.seq[17][1] ),
    .S(_0947_),
    .X(_0196_));
 sg13g2_mux2_1 _2201_ (.A0(net23),
    .A1(\simon1.seq[10][0] ),
    .S(_0950_),
    .X(_0197_));
 sg13g2_mux2_1 _2202_ (.A0(net29),
    .A1(\simon1.seq[16][1] ),
    .S(_0948_),
    .X(_0198_));
 sg13g2_mux2_1 _2203_ (.A0(net24),
    .A1(\simon1.seq[20][0] ),
    .S(_0993_),
    .X(_0199_));
 sg13g2_mux2_1 _2204_ (.A0(net31),
    .A1(\simon1.seq[1][1] ),
    .S(_0943_),
    .X(_0200_));
 sg13g2_mux2_1 _2205_ (.A0(net28),
    .A1(\simon1.seq[15][1] ),
    .S(_0949_),
    .X(_0201_));
 sg13g2_mux2_1 _2206_ (.A0(net31),
    .A1(\simon1.seq[29][1] ),
    .S(_0926_),
    .X(_0202_));
 sg13g2_and2_1 _2207_ (.A(\simon1.seq[0][1] ),
    .B(_0878_),
    .X(_0994_));
 sg13g2_a21oi_1 _2208_ (.A1(\simon1.next_random[1] ),
    .A2(_0887_),
    .Y(_0995_),
    .B1(_0994_));
 sg13g2_nand2_1 _2209_ (.Y(_0996_),
    .A(\simon1.seq[0][1] ),
    .B(_0886_));
 sg13g2_o21ai_1 _2210_ (.B1(_0996_),
    .Y(_0203_),
    .A1(net75),
    .A2(_0995_));
 sg13g2_inv_1 _2211_ (.Y(_0997_),
    .A(_0016_));
 sg13g2_nand2b_1 _2212_ (.Y(_0998_),
    .B(net83),
    .A_N(\simon1.score_rst ));
 sg13g2_buf_1 fanout32 (.A(_0892_),
    .X(net32));
 sg13g2_nor2_1 _2214_ (.A(_0997_),
    .B(_0998_),
    .Y(_0081_));
 sg13g2_xnor2_1 _2215_ (.Y(_1000_),
    .A(\simon1.score1.ones[0] ),
    .B(\simon1.score1.inc ));
 sg13g2_nor2_1 _2216_ (.A(net46),
    .B(_1000_),
    .Y(_0090_));
 sg13g2_nand2_2 _2217_ (.Y(_1001_),
    .A(\simon1.score1.ones[0] ),
    .B(\simon1.score1.inc ));
 sg13g2_nor2_1 _2218_ (.A(\simon1.score1.ones[2] ),
    .B(_0844_),
    .Y(_1002_));
 sg13g2_nor3_1 _2219_ (.A(\simon1.score1.ones[1] ),
    .B(_1001_),
    .C(_1002_),
    .Y(_1003_));
 sg13g2_a21oi_1 _2220_ (.A1(\simon1.score1.ones[1] ),
    .A2(_1001_),
    .Y(_1004_),
    .B1(_1003_));
 sg13g2_nor2_1 _2221_ (.A(net46),
    .B(_1004_),
    .Y(_0091_));
 sg13g2_nand3_1 _2222_ (.B(\simon1.score1.ones[1] ),
    .C(\simon1.score1.inc ),
    .A(\simon1.score1.ones[0] ),
    .Y(_1005_));
 sg13g2_xnor2_1 _2223_ (.Y(_1006_),
    .A(_0835_),
    .B(_1005_));
 sg13g2_nor2_1 _2224_ (.A(net46),
    .B(_1006_),
    .Y(_0092_));
 sg13g2_nor2_1 _2225_ (.A(\simon1.score1.ones[1] ),
    .B(_0835_),
    .Y(_1007_));
 sg13g2_o21ai_1 _2226_ (.B1(\simon1.score1.ones[3] ),
    .Y(_1008_),
    .A1(_1001_),
    .A2(_1007_));
 sg13g2_nor3_1 _2227_ (.A(_0835_),
    .B(\simon1.score1.ones[3] ),
    .C(_1001_),
    .Y(_1009_));
 sg13g2_o21ai_1 _2228_ (.B1(\simon1.score1.ones[1] ),
    .Y(_1010_),
    .A1(_1002_),
    .A2(_1009_));
 sg13g2_a21oi_1 _2229_ (.A1(_1008_),
    .A2(_1010_),
    .Y(_0093_),
    .B1(net46));
 sg13g2_nor4_2 _2230_ (.A(\simon1.score1.ones[1] ),
    .B(\simon1.score1.ones[2] ),
    .C(_0844_),
    .Y(_1011_),
    .D(_1001_));
 sg13g2_xnor2_1 _2231_ (.Y(_1012_),
    .A(\simon1.score1.tens[0] ),
    .B(_1011_));
 sg13g2_nor2_1 _2232_ (.A(net46),
    .B(_1012_),
    .Y(_0094_));
 sg13g2_nand2_1 _2233_ (.Y(_1013_),
    .A(\simon1.score1.tens[0] ),
    .B(_1011_));
 sg13g2_nor2b_1 _2234_ (.A(\simon1.score1.tens[2] ),
    .B_N(\simon1.score1.tens[3] ),
    .Y(_1014_));
 sg13g2_nor3_1 _2235_ (.A(\simon1.score1.tens[1] ),
    .B(_1013_),
    .C(_1014_),
    .Y(_1015_));
 sg13g2_a21oi_1 _2236_ (.A1(\simon1.score1.tens[1] ),
    .A2(_1013_),
    .Y(_1016_),
    .B1(_1015_));
 sg13g2_nor2_1 _2237_ (.A(net46),
    .B(_1016_),
    .Y(_0095_));
 sg13g2_inv_1 _2238_ (.Y(_1017_),
    .A(\simon1.score1.tens[2] ));
 sg13g2_nand3_1 _2239_ (.B(\simon1.score1.tens[1] ),
    .C(_1011_),
    .A(\simon1.score1.tens[0] ),
    .Y(_1018_));
 sg13g2_xnor2_1 _2240_ (.Y(_1019_),
    .A(_1017_),
    .B(_1018_));
 sg13g2_nor2_1 _2241_ (.A(net46),
    .B(_1019_),
    .Y(_0096_));
 sg13g2_nor2_1 _2242_ (.A(\simon1.score1.tens[1] ),
    .B(_1017_),
    .Y(_1020_));
 sg13g2_o21ai_1 _2243_ (.B1(\simon1.score1.tens[3] ),
    .Y(_1021_),
    .A1(_1013_),
    .A2(_1020_));
 sg13g2_nor3_1 _2244_ (.A(_1017_),
    .B(\simon1.score1.tens[3] ),
    .C(_1013_),
    .Y(_1022_));
 sg13g2_o21ai_1 _2245_ (.B1(\simon1.score1.tens[1] ),
    .Y(_1023_),
    .A1(_1014_),
    .A2(_1022_));
 sg13g2_a21oi_1 _2246_ (.A1(_1021_),
    .A2(_1023_),
    .Y(_0097_),
    .B1(net46));
 sg13g2_inv_1 _2247_ (.Y(_1024_),
    .A(\simon1.play1.tick_counter[30] ));
 sg13g2_or4_1 _2248_ (.A(\simon1.play1.tick_counter[22] ),
    .B(\simon1.play1.tick_counter[21] ),
    .C(\simon1.play1.tick_counter[20] ),
    .D(\simon1.play1.tick_counter[19] ),
    .X(_1025_));
 sg13g2_or2_1 _2249_ (.X(_1026_),
    .B(_1025_),
    .A(\simon1.play1.tick_counter[23] ));
 sg13g2_nor4_2 _2250_ (.A(\simon1.play1.tick_counter[26] ),
    .B(\simon1.play1.tick_counter[25] ),
    .C(\simon1.play1.tick_counter[24] ),
    .Y(_1027_),
    .D(_1026_));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31));
 sg13g2_nor3_1 _2252_ (.A(\simon1.play1.tick_counter[29] ),
    .B(\simon1.play1.tick_counter[28] ),
    .C(\simon1.play1.tick_counter[27] ),
    .Y(_1029_));
 sg13g2_and3_1 _2253_ (.X(_1030_),
    .A(_1024_),
    .B(_1027_),
    .C(_1029_));
 sg13g2_buf_1 fanout30 (.A(net32),
    .X(net30));
 sg13g2_nor4_1 _2255_ (.A(\simon1.play1.tick_counter[31] ),
    .B(\simon1.play1.tick_counter[18] ),
    .C(\simon1.play1.tick_counter[17] ),
    .D(\simon1.play1.tick_counter[16] ),
    .Y(_1032_));
 sg13g2_buf_2 fanout29 (.A(net30),
    .X(net29));
 sg13g2_buf_2 fanout28 (.A(net30),
    .X(net28));
 sg13g2_buf_1 fanout27 (.A(_0910_),
    .X(net27));
 sg13g2_buf_1 fanout26 (.A(_0910_),
    .X(net26));
 sg13g2_or3_1 _2260_ (.A(\simon1.play1.tick_counter[12] ),
    .B(\simon1.play1.tick_counter[11] ),
    .C(\simon1.play1.tick_counter[10] ),
    .X(_1037_));
 sg13g2_nand2_1 _2261_ (.Y(_1038_),
    .A(\simon1.play1.tick_counter[14] ),
    .B(\simon1.play1.tick_counter[13] ));
 sg13g2_nor4_1 _2262_ (.A(\simon1.play1.tick_counter[15] ),
    .B(\simon1.play1.tick_counter[9] ),
    .C(_1037_),
    .D(_1038_),
    .Y(_1039_));
 sg13g2_buf_1 fanout25 (.A(_0910_),
    .X(net25));
 sg13g2_nor3_1 _2264_ (.A(\simon1.play1.tick_counter[0] ),
    .B(\simon1.play1.tick_counter[1] ),
    .C(\simon1.play1.tick_counter[6] ),
    .Y(_1041_));
 sg13g2_buf_2 fanout24 (.A(net25),
    .X(net24));
 sg13g2_inv_1 _2266_ (.Y(_1043_),
    .A(\simon1.play1.tick_counter[3] ));
 sg13g2_buf_2 fanout23 (.A(net25),
    .X(net23));
 sg13g2_buf_2 fanout22 (.A(_0400_),
    .X(net22));
 sg13g2_nand2_1 _2269_ (.Y(_1046_),
    .A(\simon1.play1.tick_counter[7] ),
    .B(\simon1.play1.tick_counter[8] ));
 sg13g2_buf_2 fanout21 (.A(_0424_),
    .X(net21));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_nand2b_1 _2272_ (.Y(_1049_),
    .B(\simon1.play1.tick_counter[5] ),
    .A_N(\simon1.play1.tick_counter[4] ));
 sg13g2_nor4_1 _2273_ (.A(_1043_),
    .B(\simon1.play1.tick_counter[2] ),
    .C(_1046_),
    .D(_1049_),
    .Y(_1050_));
 sg13g2_nand3_1 _2274_ (.B(_1041_),
    .C(_1050_),
    .A(_1039_),
    .Y(_1051_));
 sg13g2_inv_1 _2275_ (.Y(_1052_),
    .A(\simon1.play1.tick_counter[14] ));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_nor2_1 _2277_ (.A(_1052_),
    .B(_0034_),
    .Y(_1054_));
 sg13g2_inv_1 _2278_ (.Y(_1055_),
    .A(\simon1.play1.tick_counter[6] ));
 sg13g2_o21ai_1 _2279_ (.B1(\simon1.play1.tick_counter[5] ),
    .Y(_1056_),
    .A1(\simon1.play1.tick_counter[3] ),
    .A2(\simon1.play1.tick_counter[4] ));
 sg13g2_a21oi_1 _2280_ (.A1(_1055_),
    .A2(_1056_),
    .Y(_1057_),
    .B1(_1046_));
 sg13g2_nand2b_1 _2281_ (.Y(_1058_),
    .B(_1039_),
    .A_N(_1057_));
 sg13g2_o21ai_1 _2282_ (.B1(_1058_),
    .Y(_1059_),
    .A1(\simon1.play1.tick_counter[15] ),
    .A2(_1054_));
 sg13g2_and4_1 _2283_ (.A(_1030_),
    .B(_1032_),
    .C(_1051_),
    .D(_1059_),
    .X(_1060_));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_nand2_1 _2285_ (.Y(_1062_),
    .A(net18),
    .B(net38));
 sg13g2_inv_1 _2286_ (.Y(_1063_),
    .A(net38));
 sg13g2_nand2_1 _2287_ (.Y(_1064_),
    .A(_0013_),
    .B(_1063_));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_nor2_1 _2290_ (.A(\simon1.play1.freq[5] ),
    .B(\simon1.play1.freq[4] ),
    .Y(_1067_));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_nor2_1 _2292_ (.A(\simon1.play1.freq[9] ),
    .B(\simon1.play1.freq[8] ),
    .Y(_1069_));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_nor2_1 _2294_ (.A(\simon1.play1.freq[7] ),
    .B(net62),
    .Y(_1071_));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_nor4_1 _2297_ (.A(\simon1.play1.freq[1] ),
    .B(\simon1.play1.freq[0] ),
    .C(net63),
    .D(\simon1.play1.freq[2] ),
    .Y(_1074_));
 sg13g2_nand4_1 _2298_ (.B(_1069_),
    .C(_1071_),
    .A(_1067_),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_nand2_1 _2300_ (.Y(_1077_),
    .A(net81),
    .B(net44));
 sg13g2_a21oi_1 _2301_ (.A1(_1062_),
    .A2(_1064_),
    .Y(_0130_),
    .B1(_1077_));
 sg13g2_nor4_1 _2302_ (.A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[9] ),
    .C(\simon1.tick_counter[11] ),
    .D(\simon1.tick_counter[10] ),
    .Y(_1078_));
 sg13g2_nor4_1 _2303_ (.A(\simon1.tick_counter[13] ),
    .B(\simon1.tick_counter[12] ),
    .C(\simon1.tick_counter[15] ),
    .D(\simon1.tick_counter[14] ),
    .Y(_1079_));
 sg13g2_nor4_1 _2304_ (.A(\simon1.tick_counter[3] ),
    .B(\simon1.tick_counter[2] ),
    .C(\simon1.tick_counter[7] ),
    .D(\simon1.tick_counter[6] ),
    .Y(_1080_));
 sg13g2_inv_1 _2305_ (.Y(_1081_),
    .A(\simon1.tick_counter[0] ));
 sg13g2_nand2_1 _2306_ (.Y(_1082_),
    .A(\simon1.tick_counter[5] ),
    .B(\simon1.tick_counter[4] ));
 sg13g2_nor3_1 _2307_ (.A(_1081_),
    .B(\simon1.tick_counter[8] ),
    .C(_1082_),
    .Y(_1083_));
 sg13g2_and4_2 _2308_ (.A(_1078_),
    .B(_1079_),
    .C(_1080_),
    .D(_1083_),
    .X(_1084_));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_inv_1 _2310_ (.Y(_1086_),
    .A(_1084_));
 sg13g2_and3_1 _2311_ (.X(_0161_),
    .A(net83),
    .B(_0036_),
    .C(_1086_));
 sg13g2_nand2_1 _2312_ (.Y(_1087_),
    .A(net83),
    .B(_1086_));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_xnor2_1 _2314_ (.Y(_1089_),
    .A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[0] ));
 sg13g2_nor2_1 _2315_ (.A(net37),
    .B(_1089_),
    .Y(_0162_));
 sg13g2_nand2_1 _2316_ (.Y(_1090_),
    .A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[0] ));
 sg13g2_xor2_1 _2317_ (.B(_1090_),
    .A(\simon1.tick_counter[2] ),
    .X(_1091_));
 sg13g2_nor2_1 _2318_ (.A(net37),
    .B(_1091_),
    .Y(_0163_));
 sg13g2_nand3_1 _2319_ (.B(\simon1.tick_counter[0] ),
    .C(\simon1.tick_counter[2] ),
    .A(\simon1.tick_counter[1] ),
    .Y(_1092_));
 sg13g2_xor2_1 _2320_ (.B(_1092_),
    .A(\simon1.tick_counter[3] ),
    .X(_1093_));
 sg13g2_nor2_1 _2321_ (.A(net37),
    .B(_1093_),
    .Y(_0164_));
 sg13g2_inv_1 _2322_ (.Y(_1094_),
    .A(\simon1.tick_counter[4] ));
 sg13g2_nand4_1 _2323_ (.B(\simon1.tick_counter[0] ),
    .C(\simon1.tick_counter[3] ),
    .A(\simon1.tick_counter[1] ),
    .Y(_1095_),
    .D(\simon1.tick_counter[2] ));
 sg13g2_xnor2_1 _2324_ (.Y(_1096_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_nor2_1 _2325_ (.A(net37),
    .B(_1096_),
    .Y(_0165_));
 sg13g2_nor2_1 _2326_ (.A(_1094_),
    .B(_1095_),
    .Y(_1097_));
 sg13g2_xnor2_1 _2327_ (.Y(_1098_),
    .A(\simon1.tick_counter[5] ),
    .B(_1097_));
 sg13g2_nor2_1 _2328_ (.A(net37),
    .B(_1098_),
    .Y(_0166_));
 sg13g2_nor2_1 _2329_ (.A(_1082_),
    .B(_1095_),
    .Y(_1099_));
 sg13g2_xnor2_1 _2330_ (.Y(_1100_),
    .A(\simon1.tick_counter[6] ),
    .B(_1099_));
 sg13g2_nor2_1 _2331_ (.A(net37),
    .B(_1100_),
    .Y(_0167_));
 sg13g2_nand2_1 _2332_ (.Y(_1101_),
    .A(\simon1.tick_counter[6] ),
    .B(_1099_));
 sg13g2_xor2_1 _2333_ (.B(_1101_),
    .A(\simon1.tick_counter[7] ),
    .X(_1102_));
 sg13g2_nor2_1 _2334_ (.A(net37),
    .B(_1102_),
    .Y(_0168_));
 sg13g2_and3_1 _2335_ (.X(_1103_),
    .A(\simon1.tick_counter[7] ),
    .B(\simon1.tick_counter[6] ),
    .C(_1099_));
 sg13g2_xnor2_1 _2336_ (.Y(_1104_),
    .A(\simon1.tick_counter[8] ),
    .B(_1103_));
 sg13g2_nor2_1 _2337_ (.A(net36),
    .B(_1104_),
    .Y(_0169_));
 sg13g2_inv_1 _2338_ (.Y(_1105_),
    .A(\simon1.tick_counter[9] ));
 sg13g2_nand2_1 _2339_ (.Y(_1106_),
    .A(\simon1.tick_counter[8] ),
    .B(_1103_));
 sg13g2_xnor2_1 _2340_ (.Y(_1107_),
    .A(_1105_),
    .B(_1106_));
 sg13g2_nor2_1 _2341_ (.A(net36),
    .B(_1107_),
    .Y(_0170_));
 sg13g2_nor2_1 _2342_ (.A(_1105_),
    .B(_1106_),
    .Y(_1108_));
 sg13g2_xnor2_1 _2343_ (.Y(_1109_),
    .A(\simon1.tick_counter[10] ),
    .B(_1108_));
 sg13g2_nor2_1 _2344_ (.A(net36),
    .B(_1109_),
    .Y(_0171_));
 sg13g2_nand2_1 _2345_ (.Y(_1110_),
    .A(\simon1.tick_counter[10] ),
    .B(_1108_));
 sg13g2_xor2_1 _2346_ (.B(_1110_),
    .A(\simon1.tick_counter[11] ),
    .X(_1111_));
 sg13g2_nor2_1 _2347_ (.A(net36),
    .B(_1111_),
    .Y(_0172_));
 sg13g2_inv_1 _2348_ (.Y(_1112_),
    .A(\simon1.tick_counter[12] ));
 sg13g2_nand3_1 _2349_ (.B(\simon1.tick_counter[10] ),
    .C(_1108_),
    .A(\simon1.tick_counter[11] ),
    .Y(_1113_));
 sg13g2_xnor2_1 _2350_ (.Y(_1114_),
    .A(_1112_),
    .B(_1113_));
 sg13g2_nor2_1 _2351_ (.A(net36),
    .B(_1114_),
    .Y(_0173_));
 sg13g2_nor2_1 _2352_ (.A(_1112_),
    .B(_1113_),
    .Y(_1115_));
 sg13g2_xnor2_1 _2353_ (.Y(_1116_),
    .A(\simon1.tick_counter[13] ),
    .B(_1115_));
 sg13g2_nor2_1 _2354_ (.A(net36),
    .B(_1116_),
    .Y(_0174_));
 sg13g2_nand2_1 _2355_ (.Y(_1117_),
    .A(\simon1.tick_counter[13] ),
    .B(_1115_));
 sg13g2_xor2_1 _2356_ (.B(_1117_),
    .A(\simon1.tick_counter[14] ),
    .X(_1118_));
 sg13g2_nor2_1 _2357_ (.A(net36),
    .B(_1118_),
    .Y(_0175_));
 sg13g2_nand3_1 _2358_ (.B(\simon1.tick_counter[14] ),
    .C(_1115_),
    .A(\simon1.tick_counter[13] ),
    .Y(_1119_));
 sg13g2_xor2_1 _2359_ (.B(_1119_),
    .A(\simon1.tick_counter[15] ),
    .X(_1120_));
 sg13g2_nor2_1 _2360_ (.A(net36),
    .B(_1120_),
    .Y(_0176_));
 sg13g2_nor2b_1 _2361_ (.A(_0763_),
    .B_N(_0875_),
    .Y(_1121_));
 sg13g2_and2_1 _2362_ (.A(_0787_),
    .B(_1121_),
    .X(_1122_));
 sg13g2_nand2b_1 _2363_ (.Y(_1123_),
    .B(net55),
    .A_N(net35));
 sg13g2_inv_1 _2364_ (.Y(_1124_),
    .A(_0032_));
 sg13g2_nand4_1 _2365_ (.B(_0739_),
    .C(net40),
    .A(_1124_),
    .Y(_1125_),
    .D(net39));
 sg13g2_nand3_1 _2366_ (.B(_1123_),
    .C(_1125_),
    .A(_1122_),
    .Y(_1126_));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_inv_1 _2368_ (.Y(_1128_),
    .A(net39));
 sg13g2_a21oi_1 _2369_ (.A1(net54),
    .A2(_1128_),
    .Y(_1129_),
    .B1(net55));
 sg13g2_nor4_1 _2370_ (.A(\simon1.seq_counter[0] ),
    .B(net76),
    .C(_1126_),
    .D(_1129_),
    .Y(_1130_));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_nand3_1 _2372_ (.B(net84),
    .C(_1126_),
    .A(\simon1.seq_counter[0] ),
    .Y(_1132_));
 sg13g2_nand2b_1 _2373_ (.Y(_0082_),
    .B(_1132_),
    .A_N(_1130_));
 sg13g2_a21oi_1 _2374_ (.A1(net55),
    .A2(_1124_),
    .Y(_1133_),
    .B1(net54));
 sg13g2_a21oi_2 _2375_ (.B1(_1133_),
    .Y(_1134_),
    .A2(net39),
    .A1(_0032_));
 sg13g2_a21oi_1 _2376_ (.A1(_0808_),
    .A2(_1134_),
    .Y(_1135_),
    .B1(_1126_));
 sg13g2_nand2_1 _2377_ (.Y(_1136_),
    .A(\simon1.seq_counter[1] ),
    .B(net82));
 sg13g2_inv_1 _2378_ (.Y(_1137_),
    .A(\simon1.seq_counter[1] ));
 sg13g2_and4_1 _2379_ (.A(_1122_),
    .B(_1123_),
    .C(_1125_),
    .D(_1134_),
    .X(_1138_));
 sg13g2_nand4_1 _2380_ (.B(_1137_),
    .C(net82),
    .A(\simon1.seq_counter[0] ),
    .Y(_1139_),
    .D(_1138_));
 sg13g2_o21ai_1 _2381_ (.B1(_1139_),
    .Y(_0083_),
    .A1(_1135_),
    .A2(_1136_));
 sg13g2_a21oi_1 _2382_ (.A1(_0791_),
    .A2(_1134_),
    .Y(_1140_),
    .B1(_1126_));
 sg13g2_nand2_1 _2383_ (.Y(_1141_),
    .A(\simon1.seq_counter[2] ),
    .B(net82));
 sg13g2_nor3_1 _2384_ (.A(\simon1.seq_counter[2] ),
    .B(net75),
    .C(_0791_),
    .Y(_1142_));
 sg13g2_nand2_1 _2385_ (.Y(_1143_),
    .A(_1138_),
    .B(_1142_));
 sg13g2_o21ai_1 _2386_ (.B1(_1143_),
    .Y(_0084_),
    .A1(_1140_),
    .A2(_1141_));
 sg13g2_nor2b_1 _2387_ (.A(_0795_),
    .B_N(_1134_),
    .Y(_1144_));
 sg13g2_nor2_1 _2388_ (.A(_1126_),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_nand2_1 _2389_ (.Y(_0211_),
    .A(\simon1.seq_counter[3] ),
    .B(net82));
 sg13g2_nand4_1 _2390_ (.B(net82),
    .C(_0795_),
    .A(_0794_),
    .Y(_0212_),
    .D(_1138_));
 sg13g2_o21ai_1 _2391_ (.B1(_0212_),
    .Y(_0085_),
    .A1(_1145_),
    .A2(_0211_));
 sg13g2_nor2b_1 _2392_ (.A(_0802_),
    .B_N(_1134_),
    .Y(_0213_));
 sg13g2_o21ai_1 _2393_ (.B1(\simon1.seq_counter[4] ),
    .Y(_0214_),
    .A1(_1126_),
    .A2(_0213_));
 sg13g2_nor2b_1 _2394_ (.A(\simon1.seq_counter[4] ),
    .B_N(_0802_),
    .Y(_0215_));
 sg13g2_nand3b_1 _2395_ (.B(_1134_),
    .C(_0215_),
    .Y(_0216_),
    .A_N(_1126_));
 sg13g2_a21oi_1 _2396_ (.A1(_0214_),
    .A2(_0216_),
    .Y(_0086_),
    .B1(net75));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[4]));
 sg13g2_xnor2_1 _2398_ (.Y(_0218_),
    .A(\simon1.play1.tick_counter[0] ),
    .B(\simon1.play1.freq[0] ));
 sg13g2_nor2_1 _2399_ (.A(net77),
    .B(_0218_),
    .Y(_0098_));
 sg13g2_nand2_1 _2400_ (.Y(_0219_),
    .A(\simon1.play1.tick_counter[0] ),
    .B(\simon1.play1.freq[0] ));
 sg13g2_xnor2_1 _2401_ (.Y(_0220_),
    .A(\simon1.play1.tick_counter[1] ),
    .B(\simon1.play1.freq[1] ));
 sg13g2_xnor2_1 _2402_ (.Y(_0221_),
    .A(_0219_),
    .B(_0220_));
 sg13g2_nor2_1 _2403_ (.A(net77),
    .B(_0221_),
    .Y(_0099_));
 sg13g2_nand2_1 _2404_ (.Y(_0222_),
    .A(\simon1.play1.tick_counter[1] ),
    .B(\simon1.play1.freq[1] ));
 sg13g2_nor2_1 _2405_ (.A(\simon1.play1.tick_counter[1] ),
    .B(\simon1.play1.freq[1] ),
    .Y(_0223_));
 sg13g2_a21o_1 _2406_ (.A2(_0222_),
    .A1(_0219_),
    .B1(_0223_),
    .X(_0224_));
 sg13g2_xnor2_1 _2407_ (.Y(_0225_),
    .A(\simon1.play1.tick_counter[2] ),
    .B(\simon1.play1.freq[2] ));
 sg13g2_xnor2_1 _2408_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_nor2_1 _2409_ (.A(net79),
    .B(_0226_),
    .Y(_0100_));
 sg13g2_and4_1 _2410_ (.A(_1067_),
    .B(_1069_),
    .C(_1071_),
    .D(_1074_),
    .X(_0227_));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_nand2_1 _2413_ (.Y(_0230_),
    .A(\simon1.play1.tick_counter[2] ),
    .B(\simon1.play1.freq[2] ));
 sg13g2_nor2_1 _2414_ (.A(\simon1.play1.tick_counter[2] ),
    .B(\simon1.play1.freq[2] ),
    .Y(_0231_));
 sg13g2_a21oi_2 _2415_ (.B1(_0231_),
    .Y(_0232_),
    .A2(_0230_),
    .A1(_0224_));
 sg13g2_xnor2_1 _2416_ (.Y(_0233_),
    .A(net63),
    .B(_0232_));
 sg13g2_xnor2_1 _2417_ (.Y(_0234_),
    .A(_1060_),
    .B(_0233_));
 sg13g2_nor2_1 _2418_ (.A(net43),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_xnor2_1 _2419_ (.Y(_0236_),
    .A(\simon1.play1.tick_counter[3] ),
    .B(_0235_));
 sg13g2_nor2_1 _2420_ (.A(net78),
    .B(_0236_),
    .Y(_0101_));
 sg13g2_a21oi_1 _2421_ (.A1(_0219_),
    .A2(_0222_),
    .Y(_0237_),
    .B1(_0223_));
 sg13g2_xnor2_1 _2422_ (.Y(_0238_),
    .A(\simon1.play1.tick_counter[3] ),
    .B(net63));
 sg13g2_nor2_1 _2423_ (.A(_0225_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a21oi_1 _2424_ (.A1(\simon1.play1.tick_counter[2] ),
    .A2(\simon1.play1.freq[2] ),
    .Y(_0240_),
    .B1(net63));
 sg13g2_nand3_1 _2425_ (.B(net63),
    .C(\simon1.play1.freq[2] ),
    .A(\simon1.play1.tick_counter[2] ),
    .Y(_0241_));
 sg13g2_o21ai_1 _2426_ (.B1(_0241_),
    .Y(_0242_),
    .A1(_1043_),
    .A2(_0240_));
 sg13g2_a21oi_2 _2427_ (.B1(_0242_),
    .Y(_0243_),
    .A2(_0239_),
    .A1(_0237_));
 sg13g2_xnor2_1 _2428_ (.Y(_0244_),
    .A(\simon1.play1.freq[4] ),
    .B(_0243_));
 sg13g2_xnor2_1 _2429_ (.Y(_0245_),
    .A(\simon1.play1.tick_counter[3] ),
    .B(_0233_));
 sg13g2_nor2_1 _2430_ (.A(_1060_),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net91),
    .D(_0082_),
    .Q_N(_1252_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net92),
    .D(_0083_),
    .Q_N(_1251_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net93),
    .D(_0084_),
    .Q_N(_1250_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net94),
    .D(_0085_),
    .Q_N(_1249_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net95),
    .D(_0086_),
    .Q_N(_1248_),
    .Q(_0004_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi ttsimon_90 (.L_HI(net90));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 _2439_ (.A(net96),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2440_ (.A(net97),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2441_ (.A(net98),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2442_ (.A(net99),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2443_ (.A(net100),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2444_ (.A(net101),
    .X(uio_oe[6]));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 _2446_ (.A(net88),
    .X(uio_out[7]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 _2448_ (.A(net89),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \simon1.millis_counter[0]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net102),
    .D(_0151_),
    .Q_N(_1189_),
    .Q(\simon1.millis_counter[0] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[1]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net103),
    .D(_0152_),
    .Q_N(_0017_),
    .Q(\simon1.millis_counter[1] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[2]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net104),
    .D(_0153_),
    .Q_N(_0018_),
    .Q(\simon1.millis_counter[2] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[3]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net105),
    .D(_0154_),
    .Q_N(_0019_),
    .Q(\simon1.millis_counter[3] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[4]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(_0155_),
    .Q_N(_0020_),
    .Q(\simon1.millis_counter[4] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[5]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net107),
    .D(_0156_),
    .Q_N(_0021_),
    .Q(\simon1.millis_counter[5] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[6]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net108),
    .D(_0157_),
    .Q_N(_0022_),
    .Q(\simon1.millis_counter[6] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[7]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net109),
    .D(_0158_),
    .Q_N(_0023_),
    .Q(\simon1.millis_counter[7] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[8]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net110),
    .D(_0159_),
    .Q_N(_0024_),
    .Q(\simon1.millis_counter[8] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[9]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net111),
    .D(_0160_),
    .Q_N(_0025_),
    .Q(\simon1.millis_counter[9] ));
 sg13g2_dfrbp_1 \simon1.next_random[0]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net112),
    .D(_0136_),
    .Q_N(_0037_),
    .Q(\simon1.next_random[0] ));
 sg13g2_dfrbp_1 \simon1.next_random[1]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net113),
    .D(_0137_),
    .Q_N(_1201_),
    .Q(\simon1.next_random[1] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[0]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net114),
    .D(_0141_),
    .Q_N(_1199_),
    .Q(\simon1.play1.freq[0] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[1]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net115),
    .D(_0142_),
    .Q_N(_1198_),
    .Q(\simon1.play1.freq[1] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[2]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net116),
    .D(_0143_),
    .Q_N(_1197_),
    .Q(\simon1.play1.freq[2] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[3]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net117),
    .D(_0144_),
    .Q_N(_1196_),
    .Q(\simon1.play1.freq[3] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[4]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net118),
    .D(_0145_),
    .Q_N(_1195_),
    .Q(\simon1.play1.freq[4] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[5]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net119),
    .D(_0146_),
    .Q_N(_1194_),
    .Q(\simon1.play1.freq[5] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[6]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net120),
    .D(_0147_),
    .Q_N(_1193_),
    .Q(\simon1.play1.freq[6] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[7]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net121),
    .D(_0148_),
    .Q_N(_1192_),
    .Q(\simon1.play1.freq[7] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[8]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net122),
    .D(_0149_),
    .Q_N(_1191_),
    .Q(\simon1.play1.freq[8] ));
 sg13g2_dfrbp_1 \simon1.play1.freq[9]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net123),
    .D(_0150_),
    .Q_N(_1190_),
    .Q(\simon1.play1.freq[9] ));
 sg13g2_dfrbp_1 \simon1.play1.sound$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net124),
    .D(_0130_),
    .Q_N(_0013_),
    .Q(net18));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[0]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net125),
    .D(_0098_),
    .Q_N(_1236_),
    .Q(\simon1.play1.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[10]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net126),
    .D(_0108_),
    .Q_N(_1226_),
    .Q(\simon1.play1.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[11]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net127),
    .D(_0109_),
    .Q_N(_1225_),
    .Q(\simon1.play1.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[12]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net128),
    .D(_0110_),
    .Q_N(_1224_),
    .Q(\simon1.play1.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[13]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net129),
    .D(_0111_),
    .Q_N(_0034_),
    .Q(\simon1.play1.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[14]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_0112_),
    .Q_N(_1223_),
    .Q(\simon1.play1.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[15]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net131),
    .D(_0113_),
    .Q_N(_1222_),
    .Q(\simon1.play1.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[16]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net132),
    .D(_0114_),
    .Q_N(_1221_),
    .Q(\simon1.play1.tick_counter[16] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[17]$_SDFFE_PN0N_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net133),
    .D(_0115_),
    .Q_N(_1220_),
    .Q(\simon1.play1.tick_counter[17] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[18]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net134),
    .D(_0116_),
    .Q_N(_1219_),
    .Q(\simon1.play1.tick_counter[18] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[19]$_SDFFE_PN0N_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_0117_),
    .Q_N(_1218_),
    .Q(\simon1.play1.tick_counter[19] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[1]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net136),
    .D(_0099_),
    .Q_N(_1235_),
    .Q(\simon1.play1.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[20]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net137),
    .D(_0118_),
    .Q_N(_1217_),
    .Q(\simon1.play1.tick_counter[20] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[21]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net138),
    .D(_0119_),
    .Q_N(_1216_),
    .Q(\simon1.play1.tick_counter[21] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[22]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net139),
    .D(_0120_),
    .Q_N(_1215_),
    .Q(\simon1.play1.tick_counter[22] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[23]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net140),
    .D(_0121_),
    .Q_N(_1214_),
    .Q(\simon1.play1.tick_counter[23] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[24]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net141),
    .D(_0122_),
    .Q_N(_1213_),
    .Q(\simon1.play1.tick_counter[24] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[25]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net142),
    .D(_0123_),
    .Q_N(_1212_),
    .Q(\simon1.play1.tick_counter[25] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[26]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net143),
    .D(_0124_),
    .Q_N(_1211_),
    .Q(\simon1.play1.tick_counter[26] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[27]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net144),
    .D(_0125_),
    .Q_N(_1210_),
    .Q(\simon1.play1.tick_counter[27] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[28]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net145),
    .D(_0126_),
    .Q_N(_1209_),
    .Q(\simon1.play1.tick_counter[28] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[29]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net146),
    .D(_0127_),
    .Q_N(_1208_),
    .Q(\simon1.play1.tick_counter[29] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[2]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net147),
    .D(_0100_),
    .Q_N(_1234_),
    .Q(\simon1.play1.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[30]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net148),
    .D(_0128_),
    .Q_N(_1207_),
    .Q(\simon1.play1.tick_counter[30] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[31]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net149),
    .D(_0129_),
    .Q_N(_1206_),
    .Q(\simon1.play1.tick_counter[31] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[3]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net150),
    .D(_0101_),
    .Q_N(_1233_),
    .Q(\simon1.play1.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[4]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net151),
    .D(_0102_),
    .Q_N(_1232_),
    .Q(\simon1.play1.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[5]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net152),
    .D(_0103_),
    .Q_N(_1231_),
    .Q(\simon1.play1.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[6]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net153),
    .D(_0104_),
    .Q_N(_1230_),
    .Q(\simon1.play1.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[7]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net154),
    .D(_0105_),
    .Q_N(_1229_),
    .Q(\simon1.play1.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[8]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net155),
    .D(_0106_),
    .Q_N(_1228_),
    .Q(\simon1.play1.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.play1.tick_counter[9]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net156),
    .D(_0107_),
    .Q_N(_1227_),
    .Q(\simon1.play1.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.score1.active_digit$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net157),
    .D(_0081_),
    .Q_N(_0016_),
    .Q(\simon1.score1.active_digit ));
 sg13g2_dfrbp_1 \simon1.score1.ena$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net158),
    .D(_0132_),
    .Q_N(_0027_),
    .Q(\simon1.score1.ena ));
 sg13g2_dfrbp_1 \simon1.score1.inc$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net159),
    .D(_0133_),
    .Q_N(_1204_),
    .Q(\simon1.score1.inc ));
 sg13g2_dfrbp_1 \simon1.score1.ones[0]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net160),
    .D(_0090_),
    .Q_N(_1244_),
    .Q(\simon1.score1.ones[0] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[1]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net161),
    .D(_0091_),
    .Q_N(_1243_),
    .Q(\simon1.score1.ones[1] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[2]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net162),
    .D(_0092_),
    .Q_N(_1242_),
    .Q(\simon1.score1.ones[2] ));
 sg13g2_dfrbp_1 \simon1.score1.ones[3]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net163),
    .D(_0093_),
    .Q_N(_1241_),
    .Q(\simon1.score1.ones[3] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[0]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net164),
    .D(_0094_),
    .Q_N(_1240_),
    .Q(\simon1.score1.tens[0] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[1]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net165),
    .D(_0095_),
    .Q_N(_1239_),
    .Q(\simon1.score1.tens[1] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[2]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net166),
    .D(_0096_),
    .Q_N(_1238_),
    .Q(\simon1.score1.tens[2] ));
 sg13g2_dfrbp_1 \simon1.score1.tens[3]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net167),
    .D(_0097_),
    .Q_N(_1237_),
    .Q(\simon1.score1.tens[3] ));
 sg13g2_dfrbp_1 \simon1.score_rst$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net168),
    .D(_0089_),
    .Q_N(_1245_),
    .Q(\simon1.score_rst ));
 sg13g2_dfrbp_1 \simon1.seq[0][0]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net169),
    .D(_0038_),
    .Q_N(_1294_),
    .Q(\simon1.seq[0][0] ));
 sg13g2_dfrbp_1 \simon1.seq[0][1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net170),
    .D(_0203_),
    .Q_N(_1146_),
    .Q(\simon1.seq[0][1] ));
 sg13g2_dfrbp_1 \simon1.seq[10][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net171),
    .D(_0197_),
    .Q_N(_1152_),
    .Q(\simon1.seq[10][0] ));
 sg13g2_dfrbp_1 \simon1.seq[10][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net172),
    .D(_0064_),
    .Q_N(_1268_),
    .Q(\simon1.seq[10][1] ));
 sg13g2_dfrbp_1 \simon1.seq[11][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net173),
    .D(_0066_),
    .Q_N(_1266_),
    .Q(\simon1.seq[11][0] ));
 sg13g2_dfrbp_1 \simon1.seq[11][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net174),
    .D(_0054_),
    .Q_N(_1278_),
    .Q(\simon1.seq[11][1] ));
 sg13g2_dfrbp_1 \simon1.seq[12][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net175),
    .D(_0065_),
    .Q_N(_1267_),
    .Q(\simon1.seq[12][0] ));
 sg13g2_dfrbp_1 \simon1.seq[12][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net176),
    .D(_0042_),
    .Q_N(_1290_),
    .Q(\simon1.seq[12][1] ));
 sg13g2_dfrbp_1 \simon1.seq[13][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net177),
    .D(_0063_),
    .Q_N(_1269_),
    .Q(\simon1.seq[13][0] ));
 sg13g2_dfrbp_1 \simon1.seq[13][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net178),
    .D(_0041_),
    .Q_N(_1291_),
    .Q(\simon1.seq[13][1] ));
 sg13g2_dfrbp_1 \simon1.seq[14][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net179),
    .D(_0062_),
    .Q_N(_1270_),
    .Q(\simon1.seq[14][0] ));
 sg13g2_dfrbp_1 \simon1.seq[14][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net180),
    .D(_0040_),
    .Q_N(_1292_),
    .Q(\simon1.seq[14][1] ));
 sg13g2_dfrbp_1 \simon1.seq[15][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net181),
    .D(_0061_),
    .Q_N(_1271_),
    .Q(\simon1.seq[15][0] ));
 sg13g2_dfrbp_1 \simon1.seq[15][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net182),
    .D(_0201_),
    .Q_N(_1148_),
    .Q(\simon1.seq[15][1] ));
 sg13g2_dfrbp_1 \simon1.seq[16][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net183),
    .D(_0060_),
    .Q_N(_1272_),
    .Q(\simon1.seq[16][0] ));
 sg13g2_dfrbp_1 \simon1.seq[16][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net184),
    .D(_0198_),
    .Q_N(_1151_),
    .Q(\simon1.seq[16][1] ));
 sg13g2_dfrbp_1 \simon1.seq[17][0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net185),
    .D(_0059_),
    .Q_N(_1273_),
    .Q(\simon1.seq[17][0] ));
 sg13g2_dfrbp_1 \simon1.seq[17][1]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net186),
    .D(_0196_),
    .Q_N(_1153_),
    .Q(\simon1.seq[17][1] ));
 sg13g2_dfrbp_1 \simon1.seq[18][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net187),
    .D(_0058_),
    .Q_N(_1274_),
    .Q(\simon1.seq[18][0] ));
 sg13g2_dfrbp_1 \simon1.seq[18][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net188),
    .D(_0187_),
    .Q_N(_1162_),
    .Q(\simon1.seq[18][1] ));
 sg13g2_dfrbp_1 \simon1.seq[19][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net189),
    .D(_0057_),
    .Q_N(_1275_),
    .Q(\simon1.seq[19][0] ));
 sg13g2_dfrbp_1 \simon1.seq[19][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net190),
    .D(_0195_),
    .Q_N(_1154_),
    .Q(\simon1.seq[19][1] ));
 sg13g2_dfrbp_1 \simon1.seq[1][0]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net191),
    .D(_0056_),
    .Q_N(_1276_),
    .Q(\simon1.seq[1][0] ));
 sg13g2_dfrbp_1 \simon1.seq[1][1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net192),
    .D(_0200_),
    .Q_N(_1149_),
    .Q(\simon1.seq[1][1] ));
 sg13g2_dfrbp_1 \simon1.seq[20][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net193),
    .D(_0199_),
    .Q_N(_1150_),
    .Q(\simon1.seq[20][0] ));
 sg13g2_dfrbp_1 \simon1.seq[20][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net194),
    .D(_0192_),
    .Q_N(_1157_),
    .Q(\simon1.seq[20][1] ));
 sg13g2_dfrbp_1 \simon1.seq[21][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net195),
    .D(_0055_),
    .Q_N(_1277_),
    .Q(\simon1.seq[21][0] ));
 sg13g2_dfrbp_1 \simon1.seq[21][1]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net196),
    .D(_0193_),
    .Q_N(_1156_),
    .Q(\simon1.seq[21][1] ));
 sg13g2_dfrbp_1 \simon1.seq[22][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net197),
    .D(_0053_),
    .Q_N(_1279_),
    .Q(\simon1.seq[22][0] ));
 sg13g2_dfrbp_1 \simon1.seq[22][1]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net198),
    .D(_0190_),
    .Q_N(_1159_),
    .Q(\simon1.seq[22][1] ));
 sg13g2_dfrbp_1 \simon1.seq[23][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net199),
    .D(_0052_),
    .Q_N(_1280_),
    .Q(\simon1.seq[23][0] ));
 sg13g2_dfrbp_1 \simon1.seq[23][1]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net200),
    .D(_0191_),
    .Q_N(_1158_),
    .Q(\simon1.seq[23][1] ));
 sg13g2_dfrbp_1 \simon1.seq[24][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net201),
    .D(_0051_),
    .Q_N(_1281_),
    .Q(\simon1.seq[24][0] ));
 sg13g2_dfrbp_1 \simon1.seq[24][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(_0194_),
    .Q_N(_1155_),
    .Q(\simon1.seq[24][1] ));
 sg13g2_dfrbp_1 \simon1.seq[25][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net203),
    .D(_0050_),
    .Q_N(_1282_),
    .Q(\simon1.seq[25][0] ));
 sg13g2_dfrbp_1 \simon1.seq[25][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net204),
    .D(_0189_),
    .Q_N(_1160_),
    .Q(\simon1.seq[25][1] ));
 sg13g2_dfrbp_1 \simon1.seq[26][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net205),
    .D(_0049_),
    .Q_N(_1283_),
    .Q(\simon1.seq[26][0] ));
 sg13g2_dfrbp_1 \simon1.seq[26][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net206),
    .D(_0188_),
    .Q_N(_1161_),
    .Q(\simon1.seq[26][1] ));
 sg13g2_dfrbp_1 \simon1.seq[27][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net207),
    .D(_0048_),
    .Q_N(_1284_),
    .Q(\simon1.seq[27][0] ));
 sg13g2_dfrbp_1 \simon1.seq[27][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net208),
    .D(_0186_),
    .Q_N(_1163_),
    .Q(\simon1.seq[27][1] ));
 sg13g2_dfrbp_1 \simon1.seq[28][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net209),
    .D(_0047_),
    .Q_N(_1285_),
    .Q(\simon1.seq[28][0] ));
 sg13g2_dfrbp_1 \simon1.seq[28][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net210),
    .D(_0131_),
    .Q_N(_1205_),
    .Q(\simon1.seq[28][1] ));
 sg13g2_dfrbp_1 \simon1.seq[29][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net211),
    .D(_0046_),
    .Q_N(_1286_),
    .Q(\simon1.seq[29][0] ));
 sg13g2_dfrbp_1 \simon1.seq[29][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net212),
    .D(_0202_),
    .Q_N(_1147_),
    .Q(\simon1.seq[29][1] ));
 sg13g2_dfrbp_1 \simon1.seq[2][0]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net213),
    .D(_0045_),
    .Q_N(_1287_),
    .Q(\simon1.seq[2][0] ));
 sg13g2_dfrbp_1 \simon1.seq[2][1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net214),
    .D(_0088_),
    .Q_N(_1302_),
    .Q(\simon1.seq[2][1] ));
 sg13g2_dfrbp_1 \simon1.seq[30][0]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net215),
    .D(_0080_),
    .Q_N(_1253_),
    .Q(\simon1.seq[30][0] ));
 sg13g2_dfrbp_1 \simon1.seq[30][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net216),
    .D(_0087_),
    .Q_N(_1247_),
    .Q(\simon1.seq[30][1] ));
 sg13g2_dfrbp_1 \simon1.seq[31][0]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net217),
    .D(_0044_),
    .Q_N(_1288_),
    .Q(\simon1.seq[31][0] ));
 sg13g2_dfrbp_1 \simon1.seq[31][1]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net218),
    .D(_0077_),
    .Q_N(_1256_),
    .Q(\simon1.seq[31][1] ));
 sg13g2_dfrbp_1 \simon1.seq[3][0]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net219),
    .D(_0043_),
    .Q_N(_1289_),
    .Q(\simon1.seq[3][0] ));
 sg13g2_dfrbp_1 \simon1.seq[3][1]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net220),
    .D(_0078_),
    .Q_N(_1255_),
    .Q(\simon1.seq[3][1] ));
 sg13g2_dfrbp_1 \simon1.seq[4][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net221),
    .D(_0079_),
    .Q_N(_1254_),
    .Q(\simon1.seq[4][0] ));
 sg13g2_dfrbp_1 \simon1.seq[4][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net222),
    .D(_0076_),
    .Q_N(_1257_),
    .Q(\simon1.seq[4][1] ));
 sg13g2_dfrbp_1 \simon1.seq[5][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net223),
    .D(_0075_),
    .Q_N(_1258_),
    .Q(\simon1.seq[5][0] ));
 sg13g2_dfrbp_1 \simon1.seq[5][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net224),
    .D(_0071_),
    .Q_N(_1262_),
    .Q(\simon1.seq[5][1] ));
 sg13g2_dfrbp_1 \simon1.seq[6][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net225),
    .D(_0074_),
    .Q_N(_1259_),
    .Q(\simon1.seq[6][0] ));
 sg13g2_dfrbp_1 \simon1.seq[6][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net226),
    .D(_0070_),
    .Q_N(_1263_),
    .Q(\simon1.seq[6][1] ));
 sg13g2_dfrbp_1 \simon1.seq[7][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net227),
    .D(_0073_),
    .Q_N(_1260_),
    .Q(\simon1.seq[7][0] ));
 sg13g2_dfrbp_1 \simon1.seq[7][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net228),
    .D(_0069_),
    .Q_N(_1264_),
    .Q(\simon1.seq[7][1] ));
 sg13g2_dfrbp_1 \simon1.seq[8][0]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net229),
    .D(_0072_),
    .Q_N(_1261_),
    .Q(\simon1.seq[8][0] ));
 sg13g2_dfrbp_1 \simon1.seq[8][1]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net230),
    .D(_0039_),
    .Q_N(_1293_),
    .Q(\simon1.seq[8][1] ));
 sg13g2_dfrbp_1 \simon1.seq[9][0]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net231),
    .D(_0068_),
    .Q_N(_1295_),
    .Q(\simon1.seq[9][0] ));
 sg13g2_dfrbp_1 \simon1.seq[9][1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net232),
    .D(_0067_),
    .Q_N(_1265_),
    .Q(\simon1.seq[9][1] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net233),
    .D(_0082_),
    .Q_N(_1172_),
    .Q(\simon1.seq_counter[0] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net234),
    .D(_0083_),
    .Q_N(_1171_),
    .Q(\simon1.seq_counter[1] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net235),
    .D(_0084_),
    .Q_N(_1170_),
    .Q(\simon1.seq_counter[2] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net236),
    .D(_0085_),
    .Q_N(_1169_),
    .Q(\simon1.seq_counter[3] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net237),
    .D(_0086_),
    .Q_N(_1168_),
    .Q(\simon1.seq_counter[4] ));
 sg13g2_dfrbp_1 \simon1.seq_length[0]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net238),
    .D(_0177_),
    .Q_N(_1173_),
    .Q(\simon1.seq_length[0] ));
 sg13g2_dfrbp_1 \simon1.seq_length[1]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net239),
    .D(_0178_),
    .Q_N(_0028_),
    .Q(\simon1.seq_length[1] ));
 sg13g2_dfrbp_1 \simon1.seq_length[2]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net240),
    .D(_0179_),
    .Q_N(_0029_),
    .Q(\simon1.seq_length[2] ));
 sg13g2_dfrbp_1 \simon1.seq_length[3]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net241),
    .D(_0180_),
    .Q_N(_0030_),
    .Q(\simon1.seq_length[3] ));
 sg13g2_dfrbp_1 \simon1.seq_length[4]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net242),
    .D(_0181_),
    .Q_N(_0031_),
    .Q(\simon1.seq_length[4] ));
 sg13g2_dfrbp_1 \simon1.state[0]$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net243),
    .D(_0005_),
    .Q_N(_1296_),
    .Q(\simon1.state[0] ));
 sg13g2_dfrbp_1 \simon1.state[1]$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net244),
    .D(_0006_),
    .Q_N(_1297_),
    .Q(\simon1.state[1] ));
 sg13g2_dfrbp_1 \simon1.state[2]$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net245),
    .D(_0007_),
    .Q_N(_1298_),
    .Q(\simon1.state[2] ));
 sg13g2_dfrbp_1 \simon1.state[3]$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net246),
    .D(_0008_),
    .Q_N(_1299_),
    .Q(\simon1.state[3] ));
 sg13g2_dfrbp_1 \simon1.state[4]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net247),
    .D(_0009_),
    .Q_N(_1300_),
    .Q(\simon1.state[4] ));
 sg13g2_dfrbp_1 \simon1.state[5]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net248),
    .D(_0010_),
    .Q_N(_0032_),
    .Q(\simon1.state[5] ));
 sg13g2_dfrbp_1 \simon1.state[6]$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net249),
    .D(_0011_),
    .Q_N(_1301_),
    .Q(\simon1.state[6] ));
 sg13g2_dfrbp_1 \simon1.state[7]$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net250),
    .D(_0012_),
    .Q_N(_0035_),
    .Q(\simon1.state[7] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[0]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net251),
    .D(_0161_),
    .Q_N(_0036_),
    .Q(\simon1.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[10]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net252),
    .D(_0171_),
    .Q_N(_1179_),
    .Q(\simon1.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[11]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net253),
    .D(_0172_),
    .Q_N(_1178_),
    .Q(\simon1.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[12]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net254),
    .D(_0173_),
    .Q_N(_1177_),
    .Q(\simon1.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[13]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net255),
    .D(_0174_),
    .Q_N(_1176_),
    .Q(\simon1.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[14]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net256),
    .D(_0175_),
    .Q_N(_1175_),
    .Q(\simon1.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[15]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net257),
    .D(_0176_),
    .Q_N(_1174_),
    .Q(\simon1.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[1]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net258),
    .D(_0162_),
    .Q_N(_1188_),
    .Q(\simon1.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[2]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net259),
    .D(_0163_),
    .Q_N(_1187_),
    .Q(\simon1.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[3]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net260),
    .D(_0164_),
    .Q_N(_1186_),
    .Q(\simon1.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net261),
    .D(_0165_),
    .Q_N(_1185_),
    .Q(\simon1.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net262),
    .D(_0166_),
    .Q_N(_1184_),
    .Q(\simon1.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[6]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net263),
    .D(_0167_),
    .Q_N(_1183_),
    .Q(\simon1.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[7]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net264),
    .D(_0168_),
    .Q_N(_1182_),
    .Q(\simon1.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[8]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net265),
    .D(_0169_),
    .Q_N(_1181_),
    .Q(\simon1.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[9]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net266),
    .D(_0170_),
    .Q_N(_1180_),
    .Q(\simon1.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[0]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net267),
    .D(_0138_),
    .Q_N(_0026_),
    .Q(\simon1.tone_sequence_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[1]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net268),
    .D(_0139_),
    .Q_N(_1200_),
    .Q(\simon1.tone_sequence_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[2]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net269),
    .D(_0140_),
    .Q_N(_0033_),
    .Q(\simon1.tone_sequence_counter[2] ));
 sg13g2_dfrbp_1 \simon1.user_input[0]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net270),
    .D(_0134_),
    .Q_N(_1203_),
    .Q(\simon1.user_input[0] ));
 sg13g2_dfrbp_1 \simon1.user_input[1]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net271),
    .D(_0135_),
    .Q_N(_1202_),
    .Q(\simon1.user_input[1] ));
 sg13g2_dfrbp_1 \uio_out[0]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net272),
    .D(_0204_),
    .Q_N(_1303_),
    .Q(net7));
 sg13g2_dfrbp_1 \uio_out[1]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net273),
    .D(_0205_),
    .Q_N(_1304_),
    .Q(net8));
 sg13g2_dfrbp_1 \uio_out[2]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net274),
    .D(_0206_),
    .Q_N(_1305_),
    .Q(net9));
 sg13g2_dfrbp_1 \uio_out[3]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net275),
    .D(_0207_),
    .Q_N(_1306_),
    .Q(net10));
 sg13g2_dfrbp_1 \uio_out[4]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net276),
    .D(_0208_),
    .Q_N(_1307_),
    .Q(net11));
 sg13g2_dfrbp_1 \uio_out[5]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net277),
    .D(_0209_),
    .Q_N(_1308_),
    .Q(net12));
 sg13g2_dfrbp_1 \uio_out[6]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net278),
    .D(_0210_),
    .Q_N(_1309_),
    .Q(net13));
 sg13g2_dfrbp_1 \uo_out[0]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net279),
    .D(_0182_),
    .Q_N(_1167_),
    .Q(net14));
 sg13g2_dfrbp_1 \uo_out[1]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net280),
    .D(_0183_),
    .Q_N(_1166_),
    .Q(net15));
 sg13g2_dfrbp_1 \uo_out[2]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net281),
    .D(_0184_),
    .Q_N(_1165_),
    .Q(net16));
 sg13g2_dfrbp_1 \uo_out[3]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net282),
    .D(_0185_),
    .Q_N(_1164_),
    .Q(net17));
 sg13g2_dfrbp_1 \uo_out[5]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net283),
    .D(_0014_),
    .Q_N(_1310_),
    .Q(net19));
 sg13g2_dfrbp_1 \uo_out[6]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net284),
    .D(_0015_),
    .Q_N(_1246_),
    .Q(net20));
 sg13g2_tiehi \simon1.millis_counter[9]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \simon1.next_random[0]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \simon1.next_random[1]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \simon1.play1.freq[0]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \simon1.play1.freq[1]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \simon1.play1.freq[2]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \simon1.play1.freq[3]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \simon1.play1.freq[4]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \simon1.play1.freq[5]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \simon1.play1.freq[6]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \simon1.play1.freq[7]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \simon1.play1.freq[8]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \simon1.play1.freq[9]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \simon1.play1.sound$_SDFFE_PP0N__124  (.L_HI(net124));
 sg13g2_tiehi \simon1.play1.tick_counter[0]$_SDFFE_PN0N__125  (.L_HI(net125));
 sg13g2_tiehi \simon1.play1.tick_counter[10]$_SDFFE_PN0N__126  (.L_HI(net126));
 sg13g2_tiehi \simon1.play1.tick_counter[11]$_SDFFE_PN0N__127  (.L_HI(net127));
 sg13g2_tiehi \simon1.play1.tick_counter[12]$_SDFFE_PN0N__128  (.L_HI(net128));
 sg13g2_tiehi \simon1.play1.tick_counter[13]$_SDFFE_PN0N__129  (.L_HI(net129));
 sg13g2_tiehi \simon1.play1.tick_counter[14]$_SDFFE_PN0N__130  (.L_HI(net130));
 sg13g2_tiehi \simon1.play1.tick_counter[15]$_SDFFE_PN0N__131  (.L_HI(net131));
 sg13g2_tiehi \simon1.play1.tick_counter[16]$_SDFFE_PN0N__132  (.L_HI(net132));
 sg13g2_tiehi \simon1.play1.tick_counter[17]$_SDFFE_PN0N__133  (.L_HI(net133));
 sg13g2_tiehi \simon1.play1.tick_counter[18]$_SDFFE_PN0N__134  (.L_HI(net134));
 sg13g2_tiehi \simon1.play1.tick_counter[19]$_SDFFE_PN0N__135  (.L_HI(net135));
 sg13g2_tiehi \simon1.play1.tick_counter[1]$_SDFFE_PN0N__136  (.L_HI(net136));
 sg13g2_tiehi \simon1.play1.tick_counter[20]$_SDFFE_PN0N__137  (.L_HI(net137));
 sg13g2_tiehi \simon1.play1.tick_counter[21]$_SDFFE_PN0N__138  (.L_HI(net138));
 sg13g2_tiehi \simon1.play1.tick_counter[22]$_SDFFE_PN0N__139  (.L_HI(net139));
 sg13g2_tiehi \simon1.play1.tick_counter[23]$_SDFFE_PN0N__140  (.L_HI(net140));
 sg13g2_tiehi \simon1.play1.tick_counter[24]$_SDFFE_PN0N__141  (.L_HI(net141));
 sg13g2_tiehi \simon1.play1.tick_counter[25]$_SDFFE_PN0N__142  (.L_HI(net142));
 sg13g2_tiehi \simon1.play1.tick_counter[26]$_SDFFE_PN0N__143  (.L_HI(net143));
 sg13g2_tiehi \simon1.play1.tick_counter[27]$_SDFFE_PN0N__144  (.L_HI(net144));
 sg13g2_tiehi \simon1.play1.tick_counter[28]$_SDFFE_PN0N__145  (.L_HI(net145));
 sg13g2_tiehi \simon1.play1.tick_counter[29]$_SDFFE_PN0N__146  (.L_HI(net146));
 sg13g2_tiehi \simon1.play1.tick_counter[2]$_SDFFE_PN0N__147  (.L_HI(net147));
 sg13g2_tiehi \simon1.play1.tick_counter[30]$_SDFFE_PN0N__148  (.L_HI(net148));
 sg13g2_tiehi \simon1.play1.tick_counter[31]$_SDFFE_PN0N__149  (.L_HI(net149));
 sg13g2_tiehi \simon1.play1.tick_counter[3]$_SDFFE_PN0N__150  (.L_HI(net150));
 sg13g2_tiehi \simon1.play1.tick_counter[4]$_SDFFE_PN0N__151  (.L_HI(net151));
 sg13g2_tiehi \simon1.play1.tick_counter[5]$_SDFFE_PN0N__152  (.L_HI(net152));
 sg13g2_tiehi \simon1.play1.tick_counter[6]$_SDFFE_PN0N__153  (.L_HI(net153));
 sg13g2_tiehi \simon1.play1.tick_counter[7]$_SDFFE_PN0N__154  (.L_HI(net154));
 sg13g2_tiehi \simon1.play1.tick_counter[8]$_SDFFE_PN0N__155  (.L_HI(net155));
 sg13g2_tiehi \simon1.play1.tick_counter[9]$_SDFFE_PN0N__156  (.L_HI(net156));
 sg13g2_tiehi \simon1.score1.active_digit$_SDFF_PP0__157  (.L_HI(net157));
 sg13g2_tiehi \simon1.score1.ena$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \simon1.score1.inc$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \simon1.score1.ones[0]$_SDFFE_PP0P__160  (.L_HI(net160));
 sg13g2_tiehi \simon1.score1.ones[1]$_SDFFE_PP0P__161  (.L_HI(net161));
 sg13g2_tiehi \simon1.score1.ones[2]$_SDFFE_PP0P__162  (.L_HI(net162));
 sg13g2_tiehi \simon1.score1.ones[3]$_SDFFE_PP0P__163  (.L_HI(net163));
 sg13g2_tiehi \simon1.score1.tens[0]$_SDFFE_PP0P__164  (.L_HI(net164));
 sg13g2_tiehi \simon1.score1.tens[1]$_SDFFE_PP0P__165  (.L_HI(net165));
 sg13g2_tiehi \simon1.score1.tens[2]$_SDFFE_PP0P__166  (.L_HI(net166));
 sg13g2_tiehi \simon1.score1.tens[3]$_SDFFE_PP0P__167  (.L_HI(net167));
 sg13g2_tiehi \simon1.score_rst$_SDFF_PN0__168  (.L_HI(net168));
 sg13g2_tiehi \simon1.seq[0][0]$_DFFE_PP__169  (.L_HI(net169));
 sg13g2_tiehi \simon1.seq[0][1]$_DFFE_PP__170  (.L_HI(net170));
 sg13g2_tiehi \simon1.seq[10][0]$_DFFE_PP__171  (.L_HI(net171));
 sg13g2_tiehi \simon1.seq[10][1]$_DFFE_PP__172  (.L_HI(net172));
 sg13g2_tiehi \simon1.seq[11][0]$_DFFE_PP__173  (.L_HI(net173));
 sg13g2_tiehi \simon1.seq[11][1]$_DFFE_PP__174  (.L_HI(net174));
 sg13g2_tiehi \simon1.seq[12][0]$_DFFE_PP__175  (.L_HI(net175));
 sg13g2_tiehi \simon1.seq[12][1]$_DFFE_PP__176  (.L_HI(net176));
 sg13g2_tiehi \simon1.seq[13][0]$_DFFE_PP__177  (.L_HI(net177));
 sg13g2_tiehi \simon1.seq[13][1]$_DFFE_PP__178  (.L_HI(net178));
 sg13g2_tiehi \simon1.seq[14][0]$_DFFE_PP__179  (.L_HI(net179));
 sg13g2_tiehi \simon1.seq[14][1]$_DFFE_PP__180  (.L_HI(net180));
 sg13g2_tiehi \simon1.seq[15][0]$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \simon1.seq[15][1]$_DFFE_PP__182  (.L_HI(net182));
 sg13g2_tiehi \simon1.seq[16][0]$_DFFE_PP__183  (.L_HI(net183));
 sg13g2_tiehi \simon1.seq[16][1]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \simon1.seq[17][0]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \simon1.seq[17][1]$_DFFE_PP__186  (.L_HI(net186));
 sg13g2_tiehi \simon1.seq[18][0]$_DFFE_PP__187  (.L_HI(net187));
 sg13g2_tiehi \simon1.seq[18][1]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \simon1.seq[19][0]$_DFFE_PP__189  (.L_HI(net189));
 sg13g2_tiehi \simon1.seq[19][1]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \simon1.seq[1][0]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \simon1.seq[1][1]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \simon1.seq[20][0]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \simon1.seq[20][1]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \simon1.seq[21][0]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \simon1.seq[21][1]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \simon1.seq[22][0]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \simon1.seq[22][1]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \simon1.seq[23][0]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \simon1.seq[23][1]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \simon1.seq[24][0]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \simon1.seq[24][1]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \simon1.seq[25][0]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \simon1.seq[25][1]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \simon1.seq[26][0]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \simon1.seq[26][1]$_DFFE_PP__206  (.L_HI(net206));
 sg13g2_tiehi \simon1.seq[27][0]$_DFFE_PP__207  (.L_HI(net207));
 sg13g2_tiehi \simon1.seq[27][1]$_DFFE_PP__208  (.L_HI(net208));
 sg13g2_tiehi \simon1.seq[28][0]$_DFFE_PP__209  (.L_HI(net209));
 sg13g2_tiehi \simon1.seq[28][1]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \simon1.seq[29][0]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \simon1.seq[29][1]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \simon1.seq[2][0]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \simon1.seq[2][1]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \simon1.seq[30][0]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \simon1.seq[30][1]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \simon1.seq[31][0]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \simon1.seq[31][1]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \simon1.seq[3][0]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \simon1.seq[3][1]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \simon1.seq[4][0]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \simon1.seq[4][1]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \simon1.seq[5][0]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \simon1.seq[5][1]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \simon1.seq[6][0]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \simon1.seq[6][1]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \simon1.seq[7][0]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \simon1.seq[7][1]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \simon1.seq[8][0]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \simon1.seq[8][1]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \simon1.seq[9][0]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \simon1.seq[9][1]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \simon1.seq_counter[0]$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \simon1.seq_counter[1]$_SDFFE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \simon1.seq_counter[2]$_SDFFE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \simon1.seq_counter[3]$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \simon1.seq_counter[4]$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \simon1.seq_length[0]$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \simon1.seq_length[1]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \simon1.seq_length[2]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \simon1.seq_length[3]$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \simon1.seq_length[4]$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \simon1.state[0]$_DFF_P__243  (.L_HI(net243));
 sg13g2_tiehi \simon1.state[1]$_DFF_P__244  (.L_HI(net244));
 sg13g2_tiehi \simon1.state[2]$_DFF_P__245  (.L_HI(net245));
 sg13g2_tiehi \simon1.state[3]$_DFF_P__246  (.L_HI(net246));
 sg13g2_tiehi \simon1.state[4]$_DFF_P__247  (.L_HI(net247));
 sg13g2_tiehi \simon1.state[5]$_DFF_P__248  (.L_HI(net248));
 sg13g2_tiehi \simon1.state[6]$_DFF_P__249  (.L_HI(net249));
 sg13g2_tiehi \simon1.state[7]$_DFF_P__250  (.L_HI(net250));
 sg13g2_tiehi \simon1.tick_counter[0]$_SDFF_PP0__251  (.L_HI(net251));
 sg13g2_tiehi \simon1.tick_counter[10]$_SDFF_PP0__252  (.L_HI(net252));
 sg13g2_tiehi \simon1.tick_counter[11]$_SDFF_PP0__253  (.L_HI(net253));
 sg13g2_tiehi \simon1.tick_counter[12]$_SDFF_PP0__254  (.L_HI(net254));
 sg13g2_tiehi \simon1.tick_counter[13]$_SDFF_PP0__255  (.L_HI(net255));
 sg13g2_tiehi \simon1.tick_counter[14]$_SDFF_PP0__256  (.L_HI(net256));
 sg13g2_tiehi \simon1.tick_counter[15]$_SDFF_PP0__257  (.L_HI(net257));
 sg13g2_tiehi \simon1.tick_counter[1]$_SDFF_PP0__258  (.L_HI(net258));
 sg13g2_tiehi \simon1.tick_counter[2]$_SDFF_PP0__259  (.L_HI(net259));
 sg13g2_tiehi \simon1.tick_counter[3]$_SDFF_PP0__260  (.L_HI(net260));
 sg13g2_tiehi \simon1.tick_counter[4]$_SDFF_PP0__261  (.L_HI(net261));
 sg13g2_tiehi \simon1.tick_counter[5]$_SDFF_PP0__262  (.L_HI(net262));
 sg13g2_tiehi \simon1.tick_counter[6]$_SDFF_PP0__263  (.L_HI(net263));
 sg13g2_tiehi \simon1.tick_counter[7]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \simon1.tick_counter[8]$_SDFF_PP0__265  (.L_HI(net265));
 sg13g2_tiehi \simon1.tick_counter[9]$_SDFF_PP0__266  (.L_HI(net266));
 sg13g2_tiehi \simon1.tone_sequence_counter[0]$_DFFE_PP__267  (.L_HI(net267));
 sg13g2_tiehi \simon1.tone_sequence_counter[1]$_DFFE_PP__268  (.L_HI(net268));
 sg13g2_tiehi \simon1.tone_sequence_counter[2]$_DFFE_PP__269  (.L_HI(net269));
 sg13g2_tiehi \simon1.user_input[0]$_DFFE_PP__270  (.L_HI(net270));
 sg13g2_tiehi \simon1.user_input[1]$_DFFE_PP__271  (.L_HI(net271));
 sg13g2_tiehi \uio_out[0]$_DFF_P__272  (.L_HI(net272));
 sg13g2_tiehi \uio_out[1]$_DFF_P__273  (.L_HI(net273));
 sg13g2_tiehi \uio_out[2]$_DFF_P__274  (.L_HI(net274));
 sg13g2_tiehi \uio_out[3]$_DFF_P__275  (.L_HI(net275));
 sg13g2_tiehi \uio_out[4]$_DFF_P__276  (.L_HI(net276));
 sg13g2_tiehi \uio_out[5]$_DFF_P__277  (.L_HI(net277));
 sg13g2_tiehi \uio_out[6]$_DFF_P__278  (.L_HI(net278));
 sg13g2_tiehi \uo_out[0]$_SDFFE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \uo_out[1]$_SDFFE_PN0P__280  (.L_HI(net280));
 sg13g2_tiehi \uo_out[2]$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \uo_out[3]$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \uo_out[5]$_DFF_P__283  (.L_HI(net283));
 sg13g2_tiehi \uo_out[6]$_DFF_P__284  (.L_HI(net284));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_inv_4 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_16 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_buf_16 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_8 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_inv_8 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_8 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_8 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_fill_8 FILLER_0_0_0 ();
 sg13g2_fill_8 FILLER_0_0_8 ();
 sg13g2_fill_8 FILLER_0_0_16 ();
 sg13g2_fill_8 FILLER_0_0_24 ();
 sg13g2_fill_8 FILLER_0_0_32 ();
 sg13g2_fill_8 FILLER_0_0_40 ();
 sg13g2_fill_2 FILLER_0_0_48 ();
 sg13g2_fill_2 FILLER_0_0_54 ();
 sg13g2_fill_2 FILLER_0_0_82 ();
 sg13g2_fill_4 FILLER_0_0_94 ();
 sg13g2_fill_2 FILLER_0_0_102 ();
 sg13g2_fill_1 FILLER_0_0_104 ();
 sg13g2_fill_2 FILLER_0_0_109 ();
 sg13g2_fill_8 FILLER_0_0_137 ();
 sg13g2_fill_2 FILLER_0_0_145 ();
 sg13g2_fill_1 FILLER_0_0_147 ();
 sg13g2_fill_4 FILLER_0_0_174 ();
 sg13g2_fill_2 FILLER_0_0_178 ();
 sg13g2_fill_8 FILLER_0_0_206 ();
 sg13g2_fill_8 FILLER_0_0_214 ();
 sg13g2_fill_8 FILLER_0_0_222 ();
 sg13g2_fill_8 FILLER_0_0_230 ();
 sg13g2_fill_8 FILLER_0_0_238 ();
 sg13g2_fill_8 FILLER_0_0_246 ();
 sg13g2_fill_8 FILLER_0_0_254 ();
 sg13g2_fill_8 FILLER_0_0_262 ();
 sg13g2_fill_8 FILLER_0_0_270 ();
 sg13g2_fill_8 FILLER_0_0_278 ();
 sg13g2_fill_8 FILLER_0_0_286 ();
 sg13g2_fill_8 FILLER_0_0_294 ();
 sg13g2_fill_8 FILLER_0_0_302 ();
 sg13g2_fill_8 FILLER_0_0_310 ();
 sg13g2_fill_4 FILLER_0_0_318 ();
 sg13g2_fill_1 FILLER_0_0_322 ();
 sg13g2_fill_8 FILLER_0_1_0 ();
 sg13g2_fill_8 FILLER_0_1_8 ();
 sg13g2_fill_8 FILLER_0_1_16 ();
 sg13g2_fill_8 FILLER_0_1_24 ();
 sg13g2_fill_2 FILLER_0_1_36 ();
 sg13g2_fill_2 FILLER_0_1_42 ();
 sg13g2_fill_4 FILLER_0_1_54 ();
 sg13g2_fill_4 FILLER_0_1_84 ();
 sg13g2_fill_1 FILLER_0_1_88 ();
 sg13g2_fill_2 FILLER_0_1_115 ();
 sg13g2_fill_1 FILLER_0_1_117 ();
 sg13g2_fill_4 FILLER_0_1_144 ();
 sg13g2_fill_1 FILLER_0_1_148 ();
 sg13g2_fill_8 FILLER_0_1_175 ();
 sg13g2_fill_4 FILLER_0_1_183 ();
 sg13g2_fill_8 FILLER_0_1_191 ();
 sg13g2_fill_4 FILLER_0_1_199 ();
 sg13g2_fill_2 FILLER_0_1_203 ();
 sg13g2_fill_8 FILLER_0_1_209 ();
 sg13g2_fill_8 FILLER_0_1_217 ();
 sg13g2_fill_8 FILLER_0_1_225 ();
 sg13g2_fill_8 FILLER_0_1_233 ();
 sg13g2_fill_8 FILLER_0_1_241 ();
 sg13g2_fill_8 FILLER_0_1_249 ();
 sg13g2_fill_8 FILLER_0_1_257 ();
 sg13g2_fill_8 FILLER_0_1_265 ();
 sg13g2_fill_8 FILLER_0_1_273 ();
 sg13g2_fill_8 FILLER_0_1_281 ();
 sg13g2_fill_8 FILLER_0_1_289 ();
 sg13g2_fill_8 FILLER_0_1_297 ();
 sg13g2_fill_8 FILLER_0_1_305 ();
 sg13g2_fill_8 FILLER_0_1_313 ();
 sg13g2_fill_2 FILLER_0_1_321 ();
 sg13g2_fill_8 FILLER_0_2_0 ();
 sg13g2_fill_8 FILLER_0_2_8 ();
 sg13g2_fill_4 FILLER_0_2_16 ();
 sg13g2_fill_2 FILLER_0_2_30 ();
 sg13g2_fill_2 FILLER_0_2_58 ();
 sg13g2_fill_4 FILLER_0_2_70 ();
 sg13g2_fill_1 FILLER_0_2_74 ();
 sg13g2_fill_2 FILLER_0_2_80 ();
 sg13g2_fill_1 FILLER_0_2_82 ();
 sg13g2_fill_2 FILLER_0_2_93 ();
 sg13g2_fill_4 FILLER_0_2_99 ();
 sg13g2_fill_4 FILLER_0_2_113 ();
 sg13g2_fill_4 FILLER_0_2_127 ();
 sg13g2_fill_2 FILLER_0_2_131 ();
 sg13g2_fill_2 FILLER_0_2_138 ();
 sg13g2_fill_1 FILLER_0_2_140 ();
 sg13g2_fill_2 FILLER_0_2_151 ();
 sg13g2_fill_2 FILLER_0_2_157 ();
 sg13g2_fill_2 FILLER_0_2_163 ();
 sg13g2_fill_1 FILLER_0_2_165 ();
 sg13g2_fill_2 FILLER_0_2_176 ();
 sg13g2_fill_8 FILLER_0_2_188 ();
 sg13g2_fill_2 FILLER_0_2_196 ();
 sg13g2_fill_8 FILLER_0_2_224 ();
 sg13g2_fill_4 FILLER_0_2_232 ();
 sg13g2_fill_8 FILLER_0_2_262 ();
 sg13g2_fill_8 FILLER_0_2_270 ();
 sg13g2_fill_8 FILLER_0_2_278 ();
 sg13g2_fill_8 FILLER_0_2_286 ();
 sg13g2_fill_8 FILLER_0_2_294 ();
 sg13g2_fill_8 FILLER_0_2_302 ();
 sg13g2_fill_8 FILLER_0_2_310 ();
 sg13g2_fill_4 FILLER_0_2_318 ();
 sg13g2_fill_1 FILLER_0_2_322 ();
 sg13g2_fill_8 FILLER_0_3_0 ();
 sg13g2_fill_8 FILLER_0_3_8 ();
 sg13g2_fill_8 FILLER_0_3_16 ();
 sg13g2_fill_4 FILLER_0_3_24 ();
 sg13g2_fill_2 FILLER_0_3_28 ();
 sg13g2_fill_1 FILLER_0_3_30 ();
 sg13g2_fill_4 FILLER_0_3_57 ();
 sg13g2_fill_2 FILLER_0_3_61 ();
 sg13g2_fill_2 FILLER_0_3_67 ();
 sg13g2_fill_1 FILLER_0_3_69 ();
 sg13g2_fill_4 FILLER_0_3_75 ();
 sg13g2_fill_4 FILLER_0_3_83 ();
 sg13g2_fill_2 FILLER_0_3_113 ();
 sg13g2_fill_1 FILLER_0_3_115 ();
 sg13g2_fill_4 FILLER_0_3_120 ();
 sg13g2_fill_2 FILLER_0_3_128 ();
 sg13g2_fill_1 FILLER_0_3_130 ();
 sg13g2_fill_2 FILLER_0_3_135 ();
 sg13g2_fill_1 FILLER_0_3_137 ();
 sg13g2_fill_4 FILLER_0_3_164 ();
 sg13g2_fill_4 FILLER_0_3_172 ();
 sg13g2_fill_1 FILLER_0_3_176 ();
 sg13g2_fill_8 FILLER_0_3_187 ();
 sg13g2_fill_8 FILLER_0_3_195 ();
 sg13g2_fill_8 FILLER_0_3_203 ();
 sg13g2_fill_8 FILLER_0_3_211 ();
 sg13g2_fill_8 FILLER_0_3_219 ();
 sg13g2_fill_4 FILLER_0_3_227 ();
 sg13g2_fill_1 FILLER_0_3_231 ();
 sg13g2_fill_2 FILLER_0_3_258 ();
 sg13g2_fill_8 FILLER_0_3_263 ();
 sg13g2_fill_4 FILLER_0_3_271 ();
 sg13g2_fill_8 FILLER_0_3_279 ();
 sg13g2_fill_8 FILLER_0_3_287 ();
 sg13g2_fill_8 FILLER_0_3_295 ();
 sg13g2_fill_8 FILLER_0_3_303 ();
 sg13g2_fill_8 FILLER_0_3_311 ();
 sg13g2_fill_4 FILLER_0_3_319 ();
 sg13g2_fill_8 FILLER_0_4_0 ();
 sg13g2_fill_8 FILLER_0_4_8 ();
 sg13g2_fill_8 FILLER_0_4_16 ();
 sg13g2_fill_1 FILLER_0_4_24 ();
 sg13g2_fill_2 FILLER_0_4_30 ();
 sg13g2_fill_4 FILLER_0_4_42 ();
 sg13g2_fill_1 FILLER_0_4_46 ();
 sg13g2_fill_2 FILLER_0_4_68 ();
 sg13g2_fill_2 FILLER_0_4_74 ();
 sg13g2_fill_1 FILLER_0_4_76 ();
 sg13g2_fill_2 FILLER_0_4_103 ();
 sg13g2_fill_2 FILLER_0_4_126 ();
 sg13g2_fill_2 FILLER_0_4_138 ();
 sg13g2_fill_2 FILLER_0_4_166 ();
 sg13g2_fill_2 FILLER_0_4_178 ();
 sg13g2_fill_1 FILLER_0_4_180 ();
 sg13g2_fill_2 FILLER_0_4_187 ();
 sg13g2_fill_2 FILLER_0_4_195 ();
 sg13g2_fill_2 FILLER_0_4_223 ();
 sg13g2_fill_8 FILLER_0_4_229 ();
 sg13g2_fill_2 FILLER_0_4_241 ();
 sg13g2_fill_8 FILLER_0_4_247 ();
 sg13g2_fill_1 FILLER_0_4_255 ();
 sg13g2_fill_2 FILLER_0_4_268 ();
 sg13g2_fill_8 FILLER_0_4_296 ();
 sg13g2_fill_8 FILLER_0_4_304 ();
 sg13g2_fill_8 FILLER_0_4_312 ();
 sg13g2_fill_2 FILLER_0_4_320 ();
 sg13g2_fill_1 FILLER_0_4_322 ();
 sg13g2_fill_8 FILLER_0_5_0 ();
 sg13g2_fill_8 FILLER_0_5_8 ();
 sg13g2_fill_8 FILLER_0_5_16 ();
 sg13g2_fill_2 FILLER_0_5_50 ();
 sg13g2_fill_2 FILLER_0_5_73 ();
 sg13g2_fill_2 FILLER_0_5_85 ();
 sg13g2_fill_2 FILLER_0_5_92 ();
 sg13g2_fill_2 FILLER_0_5_104 ();
 sg13g2_fill_2 FILLER_0_5_132 ();
 sg13g2_fill_2 FILLER_0_5_144 ();
 sg13g2_fill_2 FILLER_0_5_150 ();
 sg13g2_fill_2 FILLER_0_5_156 ();
 sg13g2_fill_2 FILLER_0_5_168 ();
 sg13g2_fill_2 FILLER_0_5_175 ();
 sg13g2_fill_1 FILLER_0_5_177 ();
 sg13g2_fill_2 FILLER_0_5_188 ();
 sg13g2_fill_2 FILLER_0_5_216 ();
 sg13g2_fill_8 FILLER_0_5_244 ();
 sg13g2_fill_1 FILLER_0_5_252 ();
 sg13g2_fill_2 FILLER_0_5_256 ();
 sg13g2_fill_2 FILLER_0_5_262 ();
 sg13g2_fill_1 FILLER_0_5_264 ();
 sg13g2_fill_2 FILLER_0_5_268 ();
 sg13g2_fill_1 FILLER_0_5_270 ();
 sg13g2_fill_2 FILLER_0_5_276 ();
 sg13g2_fill_1 FILLER_0_5_278 ();
 sg13g2_fill_4 FILLER_0_5_284 ();
 sg13g2_fill_8 FILLER_0_5_292 ();
 sg13g2_fill_8 FILLER_0_5_300 ();
 sg13g2_fill_8 FILLER_0_5_308 ();
 sg13g2_fill_4 FILLER_0_5_316 ();
 sg13g2_fill_2 FILLER_0_5_320 ();
 sg13g2_fill_1 FILLER_0_5_322 ();
 sg13g2_fill_8 FILLER_0_6_0 ();
 sg13g2_fill_8 FILLER_0_6_8 ();
 sg13g2_fill_8 FILLER_0_6_16 ();
 sg13g2_fill_8 FILLER_0_6_24 ();
 sg13g2_fill_8 FILLER_0_6_36 ();
 sg13g2_fill_4 FILLER_0_6_54 ();
 sg13g2_fill_2 FILLER_0_6_68 ();
 sg13g2_fill_2 FILLER_0_6_96 ();
 sg13g2_fill_1 FILLER_0_6_98 ();
 sg13g2_fill_2 FILLER_0_6_109 ();
 sg13g2_fill_2 FILLER_0_6_132 ();
 sg13g2_fill_2 FILLER_0_6_138 ();
 sg13g2_fill_2 FILLER_0_6_144 ();
 sg13g2_fill_2 FILLER_0_6_172 ();
 sg13g2_fill_2 FILLER_0_6_179 ();
 sg13g2_fill_2 FILLER_0_6_191 ();
 sg13g2_fill_2 FILLER_0_6_198 ();
 sg13g2_fill_2 FILLER_0_6_204 ();
 sg13g2_fill_4 FILLER_0_6_210 ();
 sg13g2_fill_2 FILLER_0_6_224 ();
 sg13g2_fill_1 FILLER_0_6_226 ();
 sg13g2_fill_2 FILLER_0_6_232 ();
 sg13g2_fill_1 FILLER_0_6_234 ();
 sg13g2_fill_2 FILLER_0_6_240 ();
 sg13g2_fill_2 FILLER_0_6_249 ();
 sg13g2_fill_4 FILLER_0_6_256 ();
 sg13g2_fill_2 FILLER_0_6_265 ();
 sg13g2_fill_4 FILLER_0_6_272 ();
 sg13g2_fill_1 FILLER_0_6_276 ();
 sg13g2_fill_8 FILLER_0_6_303 ();
 sg13g2_fill_8 FILLER_0_6_311 ();
 sg13g2_fill_4 FILLER_0_6_319 ();
 sg13g2_fill_8 FILLER_0_7_0 ();
 sg13g2_fill_8 FILLER_0_7_8 ();
 sg13g2_fill_8 FILLER_0_7_16 ();
 sg13g2_fill_8 FILLER_0_7_24 ();
 sg13g2_fill_2 FILLER_0_7_32 ();
 sg13g2_fill_2 FILLER_0_7_38 ();
 sg13g2_fill_8 FILLER_0_7_50 ();
 sg13g2_fill_8 FILLER_0_7_58 ();
 sg13g2_fill_4 FILLER_0_7_71 ();
 sg13g2_fill_1 FILLER_0_7_75 ();
 sg13g2_fill_2 FILLER_0_7_80 ();
 sg13g2_fill_1 FILLER_0_7_82 ();
 sg13g2_fill_4 FILLER_0_7_87 ();
 sg13g2_fill_8 FILLER_0_7_95 ();
 sg13g2_fill_4 FILLER_0_7_103 ();
 sg13g2_fill_2 FILLER_0_7_133 ();
 sg13g2_fill_1 FILLER_0_7_135 ();
 sg13g2_fill_4 FILLER_0_7_146 ();
 sg13g2_fill_4 FILLER_0_7_176 ();
 sg13g2_fill_4 FILLER_0_7_206 ();
 sg13g2_fill_2 FILLER_0_7_214 ();
 sg13g2_fill_1 FILLER_0_7_216 ();
 sg13g2_fill_2 FILLER_0_7_221 ();
 sg13g2_fill_1 FILLER_0_7_223 ();
 sg13g2_fill_4 FILLER_0_7_227 ();
 sg13g2_fill_2 FILLER_0_7_236 ();
 sg13g2_fill_2 FILLER_0_7_245 ();
 sg13g2_fill_4 FILLER_0_7_252 ();
 sg13g2_fill_1 FILLER_0_7_256 ();
 sg13g2_fill_2 FILLER_0_7_263 ();
 sg13g2_fill_2 FILLER_0_7_270 ();
 sg13g2_fill_2 FILLER_0_7_280 ();
 sg13g2_fill_2 FILLER_0_7_286 ();
 sg13g2_fill_2 FILLER_0_7_296 ();
 sg13g2_fill_2 FILLER_0_7_303 ();
 sg13g2_fill_1 FILLER_0_7_305 ();
 sg13g2_fill_8 FILLER_0_7_311 ();
 sg13g2_fill_4 FILLER_0_7_319 ();
 sg13g2_fill_8 FILLER_0_8_0 ();
 sg13g2_fill_8 FILLER_0_8_8 ();
 sg13g2_fill_8 FILLER_0_8_16 ();
 sg13g2_fill_2 FILLER_0_8_24 ();
 sg13g2_fill_1 FILLER_0_8_26 ();
 sg13g2_fill_2 FILLER_0_8_53 ();
 sg13g2_fill_2 FILLER_0_8_59 ();
 sg13g2_fill_4 FILLER_0_8_65 ();
 sg13g2_fill_1 FILLER_0_8_69 ();
 sg13g2_fill_2 FILLER_0_8_75 ();
 sg13g2_fill_2 FILLER_0_8_82 ();
 sg13g2_fill_2 FILLER_0_8_110 ();
 sg13g2_fill_2 FILLER_0_8_116 ();
 sg13g2_fill_1 FILLER_0_8_118 ();
 sg13g2_fill_2 FILLER_0_8_124 ();
 sg13g2_fill_8 FILLER_0_8_130 ();
 sg13g2_fill_2 FILLER_0_8_138 ();
 sg13g2_fill_2 FILLER_0_8_150 ();
 sg13g2_fill_2 FILLER_0_8_157 ();
 sg13g2_fill_2 FILLER_0_8_163 ();
 sg13g2_fill_2 FILLER_0_8_170 ();
 sg13g2_fill_2 FILLER_0_8_182 ();
 sg13g2_fill_2 FILLER_0_8_210 ();
 sg13g2_fill_1 FILLER_0_8_212 ();
 sg13g2_fill_2 FILLER_0_8_218 ();
 sg13g2_fill_2 FILLER_0_8_227 ();
 sg13g2_fill_2 FILLER_0_8_234 ();
 sg13g2_fill_2 FILLER_0_8_240 ();
 sg13g2_fill_2 FILLER_0_8_246 ();
 sg13g2_fill_2 FILLER_0_8_260 ();
 sg13g2_fill_2 FILLER_0_8_267 ();
 sg13g2_fill_2 FILLER_0_8_273 ();
 sg13g2_fill_4 FILLER_0_8_280 ();
 sg13g2_fill_2 FILLER_0_8_284 ();
 sg13g2_fill_1 FILLER_0_8_286 ();
 sg13g2_fill_4 FILLER_0_8_290 ();
 sg13g2_fill_4 FILLER_0_8_299 ();
 sg13g2_fill_8 FILLER_0_8_308 ();
 sg13g2_fill_4 FILLER_0_8_316 ();
 sg13g2_fill_2 FILLER_0_8_320 ();
 sg13g2_fill_1 FILLER_0_8_322 ();
 sg13g2_fill_8 FILLER_0_9_0 ();
 sg13g2_fill_8 FILLER_0_9_8 ();
 sg13g2_fill_8 FILLER_0_9_16 ();
 sg13g2_fill_8 FILLER_0_9_24 ();
 sg13g2_fill_4 FILLER_0_9_42 ();
 sg13g2_fill_4 FILLER_0_9_72 ();
 sg13g2_fill_1 FILLER_0_9_76 ();
 sg13g2_fill_2 FILLER_0_9_87 ();
 sg13g2_fill_1 FILLER_0_9_89 ();
 sg13g2_fill_4 FILLER_0_9_116 ();
 sg13g2_fill_2 FILLER_0_9_146 ();
 sg13g2_fill_8 FILLER_0_9_153 ();
 sg13g2_fill_4 FILLER_0_9_169 ();
 sg13g2_fill_1 FILLER_0_9_173 ();
 sg13g2_fill_2 FILLER_0_9_184 ();
 sg13g2_fill_1 FILLER_0_9_186 ();
 sg13g2_fill_2 FILLER_0_9_191 ();
 sg13g2_fill_1 FILLER_0_9_193 ();
 sg13g2_fill_2 FILLER_0_9_198 ();
 sg13g2_fill_1 FILLER_0_9_200 ();
 sg13g2_fill_4 FILLER_0_9_205 ();
 sg13g2_fill_2 FILLER_0_9_235 ();
 sg13g2_fill_2 FILLER_0_9_241 ();
 sg13g2_fill_2 FILLER_0_9_247 ();
 sg13g2_fill_2 FILLER_0_9_253 ();
 sg13g2_fill_2 FILLER_0_9_259 ();
 sg13g2_fill_4 FILLER_0_9_266 ();
 sg13g2_fill_2 FILLER_0_9_277 ();
 sg13g2_fill_4 FILLER_0_9_284 ();
 sg13g2_fill_2 FILLER_0_9_293 ();
 sg13g2_fill_2 FILLER_0_9_321 ();
 sg13g2_fill_8 FILLER_0_10_0 ();
 sg13g2_fill_8 FILLER_0_10_8 ();
 sg13g2_fill_8 FILLER_0_10_16 ();
 sg13g2_fill_8 FILLER_0_10_24 ();
 sg13g2_fill_2 FILLER_0_10_42 ();
 sg13g2_fill_2 FILLER_0_10_70 ();
 sg13g2_fill_2 FILLER_0_10_76 ();
 sg13g2_fill_2 FILLER_0_10_88 ();
 sg13g2_fill_1 FILLER_0_10_90 ();
 sg13g2_fill_2 FILLER_0_10_95 ();
 sg13g2_fill_2 FILLER_0_10_101 ();
 sg13g2_fill_2 FILLER_0_10_107 ();
 sg13g2_fill_2 FILLER_0_10_119 ();
 sg13g2_fill_2 FILLER_0_10_125 ();
 sg13g2_fill_2 FILLER_0_10_153 ();
 sg13g2_fill_2 FILLER_0_10_161 ();
 sg13g2_fill_2 FILLER_0_10_171 ();
 sg13g2_fill_1 FILLER_0_10_173 ();
 sg13g2_fill_2 FILLER_0_10_178 ();
 sg13g2_fill_1 FILLER_0_10_180 ();
 sg13g2_fill_4 FILLER_0_10_185 ();
 sg13g2_fill_4 FILLER_0_10_215 ();
 sg13g2_fill_4 FILLER_0_10_224 ();
 sg13g2_fill_2 FILLER_0_10_233 ();
 sg13g2_fill_1 FILLER_0_10_235 ();
 sg13g2_fill_2 FILLER_0_10_244 ();
 sg13g2_fill_1 FILLER_0_10_246 ();
 sg13g2_fill_2 FILLER_0_10_252 ();
 sg13g2_fill_2 FILLER_0_10_257 ();
 sg13g2_fill_2 FILLER_0_10_264 ();
 sg13g2_fill_1 FILLER_0_10_266 ();
 sg13g2_fill_2 FILLER_0_10_274 ();
 sg13g2_fill_2 FILLER_0_10_281 ();
 sg13g2_fill_2 FILLER_0_10_290 ();
 sg13g2_fill_2 FILLER_0_10_299 ();
 sg13g2_fill_4 FILLER_0_10_305 ();
 sg13g2_fill_2 FILLER_0_10_309 ();
 sg13g2_fill_1 FILLER_0_10_311 ();
 sg13g2_fill_4 FILLER_0_10_316 ();
 sg13g2_fill_2 FILLER_0_10_320 ();
 sg13g2_fill_1 FILLER_0_10_322 ();
 sg13g2_fill_8 FILLER_0_11_0 ();
 sg13g2_fill_8 FILLER_0_11_8 ();
 sg13g2_fill_8 FILLER_0_11_16 ();
 sg13g2_fill_2 FILLER_0_11_24 ();
 sg13g2_fill_1 FILLER_0_11_26 ();
 sg13g2_fill_2 FILLER_0_11_37 ();
 sg13g2_fill_2 FILLER_0_11_43 ();
 sg13g2_fill_1 FILLER_0_11_45 ();
 sg13g2_fill_2 FILLER_0_11_50 ();
 sg13g2_fill_1 FILLER_0_11_52 ();
 sg13g2_fill_2 FILLER_0_11_74 ();
 sg13g2_fill_2 FILLER_0_11_80 ();
 sg13g2_fill_2 FILLER_0_11_87 ();
 sg13g2_fill_2 FILLER_0_11_93 ();
 sg13g2_fill_2 FILLER_0_11_100 ();
 sg13g2_fill_1 FILLER_0_11_102 ();
 sg13g2_fill_2 FILLER_0_11_107 ();
 sg13g2_fill_1 FILLER_0_11_109 ();
 sg13g2_fill_2 FILLER_0_11_120 ();
 sg13g2_fill_2 FILLER_0_11_132 ();
 sg13g2_fill_4 FILLER_0_11_139 ();
 sg13g2_fill_1 FILLER_0_11_143 ();
 sg13g2_fill_4 FILLER_0_11_149 ();
 sg13g2_fill_1 FILLER_0_11_153 ();
 sg13g2_fill_2 FILLER_0_11_160 ();
 sg13g2_fill_1 FILLER_0_11_162 ();
 sg13g2_fill_4 FILLER_0_11_168 ();
 sg13g2_fill_1 FILLER_0_11_172 ();
 sg13g2_fill_4 FILLER_0_11_177 ();
 sg13g2_fill_2 FILLER_0_11_191 ();
 sg13g2_fill_2 FILLER_0_11_219 ();
 sg13g2_fill_2 FILLER_0_11_226 ();
 sg13g2_fill_1 FILLER_0_11_228 ();
 sg13g2_fill_2 FILLER_0_11_234 ();
 sg13g2_fill_4 FILLER_0_11_244 ();
 sg13g2_fill_2 FILLER_0_11_248 ();
 sg13g2_fill_1 FILLER_0_11_250 ();
 sg13g2_fill_2 FILLER_0_11_258 ();
 sg13g2_fill_2 FILLER_0_11_265 ();
 sg13g2_fill_4 FILLER_0_11_272 ();
 sg13g2_fill_1 FILLER_0_11_276 ();
 sg13g2_fill_4 FILLER_0_11_283 ();
 sg13g2_fill_1 FILLER_0_11_287 ();
 sg13g2_fill_2 FILLER_0_11_293 ();
 sg13g2_fill_2 FILLER_0_11_321 ();
 sg13g2_fill_8 FILLER_0_12_0 ();
 sg13g2_fill_8 FILLER_0_12_8 ();
 sg13g2_fill_8 FILLER_0_12_16 ();
 sg13g2_fill_4 FILLER_0_12_24 ();
 sg13g2_fill_2 FILLER_0_12_28 ();
 sg13g2_fill_2 FILLER_0_12_34 ();
 sg13g2_fill_2 FILLER_0_12_62 ();
 sg13g2_fill_1 FILLER_0_12_64 ();
 sg13g2_fill_2 FILLER_0_12_91 ();
 sg13g2_fill_2 FILLER_0_12_97 ();
 sg13g2_fill_1 FILLER_0_12_99 ();
 sg13g2_fill_2 FILLER_0_12_104 ();
 sg13g2_fill_2 FILLER_0_12_110 ();
 sg13g2_fill_2 FILLER_0_12_116 ();
 sg13g2_fill_2 FILLER_0_12_144 ();
 sg13g2_fill_2 FILLER_0_12_151 ();
 sg13g2_fill_2 FILLER_0_12_161 ();
 sg13g2_fill_2 FILLER_0_12_167 ();
 sg13g2_fill_2 FILLER_0_12_174 ();
 sg13g2_fill_1 FILLER_0_12_176 ();
 sg13g2_fill_2 FILLER_0_12_183 ();
 sg13g2_fill_2 FILLER_0_12_190 ();
 sg13g2_fill_4 FILLER_0_12_202 ();
 sg13g2_fill_2 FILLER_0_12_216 ();
 sg13g2_fill_2 FILLER_0_12_223 ();
 sg13g2_fill_4 FILLER_0_12_230 ();
 sg13g2_fill_2 FILLER_0_12_234 ();
 sg13g2_fill_2 FILLER_0_12_261 ();
 sg13g2_fill_2 FILLER_0_12_268 ();
 sg13g2_fill_2 FILLER_0_12_275 ();
 sg13g2_fill_1 FILLER_0_12_277 ();
 sg13g2_fill_2 FILLER_0_12_284 ();
 sg13g2_fill_4 FILLER_0_12_290 ();
 sg13g2_fill_2 FILLER_0_12_294 ();
 sg13g2_fill_4 FILLER_0_12_301 ();
 sg13g2_fill_1 FILLER_0_12_305 ();
 sg13g2_fill_2 FILLER_0_12_313 ();
 sg13g2_fill_4 FILLER_0_12_319 ();
 sg13g2_fill_8 FILLER_0_13_0 ();
 sg13g2_fill_8 FILLER_0_13_8 ();
 sg13g2_fill_8 FILLER_0_13_16 ();
 sg13g2_fill_4 FILLER_0_13_24 ();
 sg13g2_fill_2 FILLER_0_13_38 ();
 sg13g2_fill_4 FILLER_0_13_44 ();
 sg13g2_fill_2 FILLER_0_13_48 ();
 sg13g2_fill_2 FILLER_0_13_71 ();
 sg13g2_fill_2 FILLER_0_13_83 ();
 sg13g2_fill_2 FILLER_0_13_93 ();
 sg13g2_fill_4 FILLER_0_13_100 ();
 sg13g2_fill_2 FILLER_0_13_104 ();
 sg13g2_fill_2 FILLER_0_13_116 ();
 sg13g2_fill_2 FILLER_0_13_144 ();
 sg13g2_fill_2 FILLER_0_13_152 ();
 sg13g2_fill_2 FILLER_0_13_160 ();
 sg13g2_fill_2 FILLER_0_13_166 ();
 sg13g2_fill_2 FILLER_0_13_173 ();
 sg13g2_fill_1 FILLER_0_13_175 ();
 sg13g2_fill_2 FILLER_0_13_181 ();
 sg13g2_fill_1 FILLER_0_13_183 ();
 sg13g2_fill_4 FILLER_0_13_190 ();
 sg13g2_fill_4 FILLER_0_13_199 ();
 sg13g2_fill_2 FILLER_0_13_207 ();
 sg13g2_fill_4 FILLER_0_13_213 ();
 sg13g2_fill_2 FILLER_0_13_217 ();
 sg13g2_fill_1 FILLER_0_13_219 ();
 sg13g2_fill_2 FILLER_0_13_246 ();
 sg13g2_fill_4 FILLER_0_13_253 ();
 sg13g2_fill_4 FILLER_0_13_262 ();
 sg13g2_fill_2 FILLER_0_13_271 ();
 sg13g2_fill_4 FILLER_0_13_279 ();
 sg13g2_fill_2 FILLER_0_13_293 ();
 sg13g2_fill_2 FILLER_0_13_321 ();
 sg13g2_fill_8 FILLER_0_14_0 ();
 sg13g2_fill_8 FILLER_0_14_8 ();
 sg13g2_fill_8 FILLER_0_14_16 ();
 sg13g2_fill_2 FILLER_0_14_24 ();
 sg13g2_fill_1 FILLER_0_14_26 ();
 sg13g2_fill_4 FILLER_0_14_53 ();
 sg13g2_fill_2 FILLER_0_14_83 ();
 sg13g2_fill_4 FILLER_0_14_91 ();
 sg13g2_fill_4 FILLER_0_14_100 ();
 sg13g2_fill_2 FILLER_0_14_104 ();
 sg13g2_fill_4 FILLER_0_14_116 ();
 sg13g2_fill_1 FILLER_0_14_120 ();
 sg13g2_fill_2 FILLER_0_14_125 ();
 sg13g2_fill_2 FILLER_0_14_137 ();
 sg13g2_fill_1 FILLER_0_14_139 ();
 sg13g2_fill_2 FILLER_0_14_145 ();
 sg13g2_fill_2 FILLER_0_14_152 ();
 sg13g2_fill_2 FILLER_0_14_162 ();
 sg13g2_fill_2 FILLER_0_14_172 ();
 sg13g2_fill_1 FILLER_0_14_174 ();
 sg13g2_fill_2 FILLER_0_14_183 ();
 sg13g2_fill_2 FILLER_0_14_193 ();
 sg13g2_fill_2 FILLER_0_14_221 ();
 sg13g2_fill_1 FILLER_0_14_223 ();
 sg13g2_fill_2 FILLER_0_14_250 ();
 sg13g2_fill_1 FILLER_0_14_252 ();
 sg13g2_fill_2 FILLER_0_14_258 ();
 sg13g2_fill_2 FILLER_0_14_264 ();
 sg13g2_fill_4 FILLER_0_14_270 ();
 sg13g2_fill_1 FILLER_0_14_274 ();
 sg13g2_fill_2 FILLER_0_14_281 ();
 sg13g2_fill_1 FILLER_0_14_283 ();
 sg13g2_fill_2 FILLER_0_14_290 ();
 sg13g2_fill_1 FILLER_0_14_292 ();
 sg13g2_fill_4 FILLER_0_14_298 ();
 sg13g2_fill_2 FILLER_0_14_306 ();
 sg13g2_fill_2 FILLER_0_14_311 ();
 sg13g2_fill_4 FILLER_0_14_318 ();
 sg13g2_fill_1 FILLER_0_14_322 ();
 sg13g2_fill_8 FILLER_0_15_0 ();
 sg13g2_fill_8 FILLER_0_15_8 ();
 sg13g2_fill_8 FILLER_0_15_16 ();
 sg13g2_fill_8 FILLER_0_15_24 ();
 sg13g2_fill_4 FILLER_0_15_36 ();
 sg13g2_fill_1 FILLER_0_15_40 ();
 sg13g2_fill_2 FILLER_0_15_45 ();
 sg13g2_fill_2 FILLER_0_15_51 ();
 sg13g2_fill_2 FILLER_0_15_63 ();
 sg13g2_fill_4 FILLER_0_15_69 ();
 sg13g2_fill_2 FILLER_0_15_73 ();
 sg13g2_fill_4 FILLER_0_15_85 ();
 sg13g2_fill_1 FILLER_0_15_89 ();
 sg13g2_fill_2 FILLER_0_15_95 ();
 sg13g2_fill_2 FILLER_0_15_102 ();
 sg13g2_fill_2 FILLER_0_15_108 ();
 sg13g2_fill_4 FILLER_0_15_114 ();
 sg13g2_fill_1 FILLER_0_15_118 ();
 sg13g2_fill_2 FILLER_0_15_145 ();
 sg13g2_fill_2 FILLER_0_15_152 ();
 sg13g2_fill_4 FILLER_0_15_159 ();
 sg13g2_fill_1 FILLER_0_15_163 ();
 sg13g2_fill_4 FILLER_0_15_170 ();
 sg13g2_fill_1 FILLER_0_15_174 ();
 sg13g2_fill_4 FILLER_0_15_181 ();
 sg13g2_fill_1 FILLER_0_15_185 ();
 sg13g2_fill_4 FILLER_0_15_192 ();
 sg13g2_fill_2 FILLER_0_15_196 ();
 sg13g2_fill_2 FILLER_0_15_202 ();
 sg13g2_fill_2 FILLER_0_15_230 ();
 sg13g2_fill_2 FILLER_0_15_236 ();
 sg13g2_fill_2 FILLER_0_15_242 ();
 sg13g2_fill_2 FILLER_0_15_248 ();
 sg13g2_fill_4 FILLER_0_15_255 ();
 sg13g2_fill_2 FILLER_0_15_264 ();
 sg13g2_fill_2 FILLER_0_15_270 ();
 sg13g2_fill_2 FILLER_0_15_276 ();
 sg13g2_fill_8 FILLER_0_15_282 ();
 sg13g2_fill_8 FILLER_0_15_290 ();
 sg13g2_fill_1 FILLER_0_15_298 ();
 sg13g2_fill_2 FILLER_0_15_305 ();
 sg13g2_fill_2 FILLER_0_15_315 ();
 sg13g2_fill_2 FILLER_0_15_321 ();
 sg13g2_fill_8 FILLER_0_16_0 ();
 sg13g2_fill_8 FILLER_0_16_8 ();
 sg13g2_fill_8 FILLER_0_16_16 ();
 sg13g2_fill_2 FILLER_0_16_34 ();
 sg13g2_fill_2 FILLER_0_16_62 ();
 sg13g2_fill_1 FILLER_0_16_64 ();
 sg13g2_fill_4 FILLER_0_16_69 ();
 sg13g2_fill_2 FILLER_0_16_73 ();
 sg13g2_fill_4 FILLER_0_16_85 ();
 sg13g2_fill_2 FILLER_0_16_89 ();
 sg13g2_fill_2 FILLER_0_16_96 ();
 sg13g2_fill_2 FILLER_0_16_101 ();
 sg13g2_fill_4 FILLER_0_16_108 ();
 sg13g2_fill_2 FILLER_0_16_122 ();
 sg13g2_fill_2 FILLER_0_16_150 ();
 sg13g2_fill_1 FILLER_0_16_152 ();
 sg13g2_fill_2 FILLER_0_16_158 ();
 sg13g2_fill_4 FILLER_0_16_166 ();
 sg13g2_fill_2 FILLER_0_16_175 ();
 sg13g2_fill_4 FILLER_0_16_181 ();
 sg13g2_fill_2 FILLER_0_16_195 ();
 sg13g2_fill_4 FILLER_0_16_207 ();
 sg13g2_fill_1 FILLER_0_16_211 ();
 sg13g2_fill_4 FILLER_0_16_238 ();
 sg13g2_fill_2 FILLER_0_16_242 ();
 sg13g2_fill_1 FILLER_0_16_244 ();
 sg13g2_fill_2 FILLER_0_16_250 ();
 sg13g2_fill_2 FILLER_0_16_257 ();
 sg13g2_fill_1 FILLER_0_16_259 ();
 sg13g2_fill_4 FILLER_0_16_264 ();
 sg13g2_fill_2 FILLER_0_16_275 ();
 sg13g2_fill_4 FILLER_0_16_282 ();
 sg13g2_fill_4 FILLER_0_16_291 ();
 sg13g2_fill_2 FILLER_0_16_321 ();
 sg13g2_fill_8 FILLER_0_17_0 ();
 sg13g2_fill_8 FILLER_0_17_8 ();
 sg13g2_fill_8 FILLER_0_17_16 ();
 sg13g2_fill_1 FILLER_0_17_24 ();
 sg13g2_fill_2 FILLER_0_17_35 ();
 sg13g2_fill_4 FILLER_0_17_63 ();
 sg13g2_fill_1 FILLER_0_17_67 ();
 sg13g2_fill_2 FILLER_0_17_73 ();
 sg13g2_fill_4 FILLER_0_17_80 ();
 sg13g2_fill_2 FILLER_0_17_84 ();
 sg13g2_fill_1 FILLER_0_17_86 ();
 sg13g2_fill_2 FILLER_0_17_92 ();
 sg13g2_fill_4 FILLER_0_17_101 ();
 sg13g2_fill_2 FILLER_0_17_105 ();
 sg13g2_fill_2 FILLER_0_17_117 ();
 sg13g2_fill_2 FILLER_0_17_144 ();
 sg13g2_fill_2 FILLER_0_17_150 ();
 sg13g2_fill_2 FILLER_0_17_157 ();
 sg13g2_fill_2 FILLER_0_17_164 ();
 sg13g2_fill_4 FILLER_0_17_170 ();
 sg13g2_fill_2 FILLER_0_17_179 ();
 sg13g2_fill_1 FILLER_0_17_181 ();
 sg13g2_fill_2 FILLER_0_17_187 ();
 sg13g2_fill_1 FILLER_0_17_189 ();
 sg13g2_fill_2 FILLER_0_17_216 ();
 sg13g2_fill_4 FILLER_0_17_222 ();
 sg13g2_fill_1 FILLER_0_17_226 ();
 sg13g2_fill_2 FILLER_0_17_235 ();
 sg13g2_fill_1 FILLER_0_17_237 ();
 sg13g2_fill_2 FILLER_0_17_244 ();
 sg13g2_fill_1 FILLER_0_17_246 ();
 sg13g2_fill_2 FILLER_0_17_273 ();
 sg13g2_fill_4 FILLER_0_17_280 ();
 sg13g2_fill_2 FILLER_0_17_284 ();
 sg13g2_fill_4 FILLER_0_17_294 ();
 sg13g2_fill_2 FILLER_0_17_302 ();
 sg13g2_fill_4 FILLER_0_17_308 ();
 sg13g2_fill_2 FILLER_0_17_312 ();
 sg13g2_fill_1 FILLER_0_17_322 ();
 sg13g2_fill_8 FILLER_0_18_0 ();
 sg13g2_fill_8 FILLER_0_18_8 ();
 sg13g2_fill_8 FILLER_0_18_16 ();
 sg13g2_fill_8 FILLER_0_18_24 ();
 sg13g2_fill_8 FILLER_0_18_32 ();
 sg13g2_fill_4 FILLER_0_18_40 ();
 sg13g2_fill_2 FILLER_0_18_44 ();
 sg13g2_fill_4 FILLER_0_18_50 ();
 sg13g2_fill_1 FILLER_0_18_54 ();
 sg13g2_fill_2 FILLER_0_18_59 ();
 sg13g2_fill_2 FILLER_0_18_65 ();
 sg13g2_fill_2 FILLER_0_18_71 ();
 sg13g2_fill_2 FILLER_0_18_78 ();
 sg13g2_fill_4 FILLER_0_18_85 ();
 sg13g2_fill_2 FILLER_0_18_89 ();
 sg13g2_fill_1 FILLER_0_18_91 ();
 sg13g2_fill_2 FILLER_0_18_99 ();
 sg13g2_fill_2 FILLER_0_18_105 ();
 sg13g2_fill_2 FILLER_0_18_111 ();
 sg13g2_fill_2 FILLER_0_18_123 ();
 sg13g2_fill_2 FILLER_0_18_151 ();
 sg13g2_fill_1 FILLER_0_18_153 ();
 sg13g2_fill_2 FILLER_0_18_160 ();
 sg13g2_fill_4 FILLER_0_18_167 ();
 sg13g2_fill_2 FILLER_0_18_171 ();
 sg13g2_fill_2 FILLER_0_18_178 ();
 sg13g2_fill_2 FILLER_0_18_190 ();
 sg13g2_fill_2 FILLER_0_18_197 ();
 sg13g2_fill_1 FILLER_0_18_199 ();
 sg13g2_fill_4 FILLER_0_18_226 ();
 sg13g2_fill_2 FILLER_0_18_230 ();
 sg13g2_fill_1 FILLER_0_18_232 ();
 sg13g2_fill_2 FILLER_0_18_238 ();
 sg13g2_fill_2 FILLER_0_18_245 ();
 sg13g2_fill_2 FILLER_0_18_251 ();
 sg13g2_fill_2 FILLER_0_18_258 ();
 sg13g2_fill_4 FILLER_0_18_264 ();
 sg13g2_fill_2 FILLER_0_18_273 ();
 sg13g2_fill_4 FILLER_0_18_279 ();
 sg13g2_fill_2 FILLER_0_18_287 ();
 sg13g2_fill_2 FILLER_0_18_292 ();
 sg13g2_fill_4 FILLER_0_18_297 ();
 sg13g2_fill_1 FILLER_0_18_301 ();
 sg13g2_fill_4 FILLER_0_18_306 ();
 sg13g2_fill_1 FILLER_0_18_310 ();
 sg13g2_fill_2 FILLER_0_18_316 ();
 sg13g2_fill_2 FILLER_0_18_321 ();
 sg13g2_fill_8 FILLER_0_19_0 ();
 sg13g2_fill_8 FILLER_0_19_8 ();
 sg13g2_fill_8 FILLER_0_19_16 ();
 sg13g2_fill_4 FILLER_0_19_24 ();
 sg13g2_fill_2 FILLER_0_19_32 ();
 sg13g2_fill_1 FILLER_0_19_34 ();
 sg13g2_fill_2 FILLER_0_19_39 ();
 sg13g2_fill_8 FILLER_0_19_45 ();
 sg13g2_fill_2 FILLER_0_19_53 ();
 sg13g2_fill_1 FILLER_0_19_55 ();
 sg13g2_fill_2 FILLER_0_19_77 ();
 sg13g2_fill_1 FILLER_0_19_79 ();
 sg13g2_fill_2 FILLER_0_19_86 ();
 sg13g2_fill_2 FILLER_0_19_93 ();
 sg13g2_fill_2 FILLER_0_19_100 ();
 sg13g2_fill_1 FILLER_0_19_102 ();
 sg13g2_fill_4 FILLER_0_19_108 ();
 sg13g2_fill_1 FILLER_0_19_112 ();
 sg13g2_fill_2 FILLER_0_19_123 ();
 sg13g2_fill_4 FILLER_0_19_151 ();
 sg13g2_fill_4 FILLER_0_19_161 ();
 sg13g2_fill_1 FILLER_0_19_165 ();
 sg13g2_fill_2 FILLER_0_19_171 ();
 sg13g2_fill_2 FILLER_0_19_177 ();
 sg13g2_fill_2 FILLER_0_19_183 ();
 sg13g2_fill_2 FILLER_0_19_189 ();
 sg13g2_fill_1 FILLER_0_19_191 ();
 sg13g2_fill_2 FILLER_0_19_202 ();
 sg13g2_fill_2 FILLER_0_19_209 ();
 sg13g2_fill_2 FILLER_0_19_216 ();
 sg13g2_fill_4 FILLER_0_19_222 ();
 sg13g2_fill_2 FILLER_0_19_231 ();
 sg13g2_fill_2 FILLER_0_19_237 ();
 sg13g2_fill_2 FILLER_0_19_244 ();
 sg13g2_fill_2 FILLER_0_19_251 ();
 sg13g2_fill_4 FILLER_0_19_279 ();
 sg13g2_fill_4 FILLER_0_19_289 ();
 sg13g2_fill_2 FILLER_0_19_300 ();
 sg13g2_fill_2 FILLER_0_19_307 ();
 sg13g2_fill_4 FILLER_0_19_319 ();
 sg13g2_fill_8 FILLER_0_20_0 ();
 sg13g2_fill_8 FILLER_0_20_8 ();
 sg13g2_fill_8 FILLER_0_20_16 ();
 sg13g2_fill_2 FILLER_0_20_34 ();
 sg13g2_fill_4 FILLER_0_20_62 ();
 sg13g2_fill_2 FILLER_0_20_66 ();
 sg13g2_fill_1 FILLER_0_20_68 ();
 sg13g2_fill_2 FILLER_0_20_95 ();
 sg13g2_fill_1 FILLER_0_20_97 ();
 sg13g2_fill_2 FILLER_0_20_102 ();
 sg13g2_fill_2 FILLER_0_20_108 ();
 sg13g2_fill_2 FILLER_0_20_114 ();
 sg13g2_fill_2 FILLER_0_20_121 ();
 sg13g2_fill_4 FILLER_0_20_149 ();
 sg13g2_fill_2 FILLER_0_20_159 ();
 sg13g2_fill_2 FILLER_0_20_166 ();
 sg13g2_fill_2 FILLER_0_20_178 ();
 sg13g2_fill_2 FILLER_0_20_184 ();
 sg13g2_fill_2 FILLER_0_20_190 ();
 sg13g2_fill_2 FILLER_0_20_202 ();
 sg13g2_fill_2 FILLER_0_20_214 ();
 sg13g2_fill_1 FILLER_0_20_216 ();
 sg13g2_fill_2 FILLER_0_20_243 ();
 sg13g2_fill_2 FILLER_0_20_255 ();
 sg13g2_fill_2 FILLER_0_20_262 ();
 sg13g2_fill_4 FILLER_0_20_270 ();
 sg13g2_fill_4 FILLER_0_20_279 ();
 sg13g2_fill_2 FILLER_0_20_291 ();
 sg13g2_fill_2 FILLER_0_20_298 ();
 sg13g2_fill_2 FILLER_0_20_305 ();
 sg13g2_fill_2 FILLER_0_20_312 ();
 sg13g2_fill_4 FILLER_0_20_319 ();
 sg13g2_fill_8 FILLER_0_21_0 ();
 sg13g2_fill_8 FILLER_0_21_8 ();
 sg13g2_fill_8 FILLER_0_21_16 ();
 sg13g2_fill_2 FILLER_0_21_34 ();
 sg13g2_fill_2 FILLER_0_21_62 ();
 sg13g2_fill_4 FILLER_0_21_74 ();
 sg13g2_fill_2 FILLER_0_21_78 ();
 sg13g2_fill_2 FILLER_0_21_84 ();
 sg13g2_fill_8 FILLER_0_21_90 ();
 sg13g2_fill_8 FILLER_0_21_98 ();
 sg13g2_fill_2 FILLER_0_21_110 ();
 sg13g2_fill_2 FILLER_0_21_122 ();
 sg13g2_fill_4 FILLER_0_21_150 ();
 sg13g2_fill_2 FILLER_0_21_154 ();
 sg13g2_fill_4 FILLER_0_21_161 ();
 sg13g2_fill_1 FILLER_0_21_165 ();
 sg13g2_fill_2 FILLER_0_21_176 ();
 sg13g2_fill_4 FILLER_0_21_204 ();
 sg13g2_fill_1 FILLER_0_21_208 ();
 sg13g2_fill_4 FILLER_0_21_219 ();
 sg13g2_fill_2 FILLER_0_21_223 ();
 sg13g2_fill_2 FILLER_0_21_230 ();
 sg13g2_fill_2 FILLER_0_21_237 ();
 sg13g2_fill_2 FILLER_0_21_243 ();
 sg13g2_fill_2 FILLER_0_21_252 ();
 sg13g2_fill_2 FILLER_0_21_260 ();
 sg13g2_fill_4 FILLER_0_21_268 ();
 sg13g2_fill_4 FILLER_0_21_280 ();
 sg13g2_fill_1 FILLER_0_21_284 ();
 sg13g2_fill_4 FILLER_0_21_289 ();
 sg13g2_fill_2 FILLER_0_21_293 ();
 sg13g2_fill_2 FILLER_0_21_321 ();
 sg13g2_fill_8 FILLER_0_22_0 ();
 sg13g2_fill_8 FILLER_0_22_8 ();
 sg13g2_fill_8 FILLER_0_22_16 ();
 sg13g2_fill_8 FILLER_0_22_24 ();
 sg13g2_fill_1 FILLER_0_22_32 ();
 sg13g2_fill_2 FILLER_0_22_43 ();
 sg13g2_fill_1 FILLER_0_22_45 ();
 sg13g2_fill_4 FILLER_0_22_50 ();
 sg13g2_fill_4 FILLER_0_22_75 ();
 sg13g2_fill_8 FILLER_0_22_105 ();
 sg13g2_fill_4 FILLER_0_22_113 ();
 sg13g2_fill_2 FILLER_0_22_127 ();
 sg13g2_fill_2 FILLER_0_22_133 ();
 sg13g2_fill_1 FILLER_0_22_135 ();
 sg13g2_fill_4 FILLER_0_22_162 ();
 sg13g2_fill_4 FILLER_0_22_171 ();
 sg13g2_fill_4 FILLER_0_22_201 ();
 sg13g2_fill_1 FILLER_0_22_205 ();
 sg13g2_fill_2 FILLER_0_22_211 ();
 sg13g2_fill_1 FILLER_0_22_213 ();
 sg13g2_fill_4 FILLER_0_22_240 ();
 sg13g2_fill_1 FILLER_0_22_244 ();
 sg13g2_fill_2 FILLER_0_22_250 ();
 sg13g2_fill_2 FILLER_0_22_257 ();
 sg13g2_fill_2 FILLER_0_22_264 ();
 sg13g2_fill_2 FILLER_0_22_271 ();
 sg13g2_fill_1 FILLER_0_22_273 ();
 sg13g2_fill_4 FILLER_0_22_280 ();
 sg13g2_fill_2 FILLER_0_22_284 ();
 sg13g2_fill_4 FILLER_0_22_290 ();
 sg13g2_fill_2 FILLER_0_22_294 ();
 sg13g2_fill_2 FILLER_0_22_300 ();
 sg13g2_fill_2 FILLER_0_22_306 ();
 sg13g2_fill_8 FILLER_0_22_312 ();
 sg13g2_fill_2 FILLER_0_22_320 ();
 sg13g2_fill_1 FILLER_0_22_322 ();
 sg13g2_fill_8 FILLER_0_23_0 ();
 sg13g2_fill_8 FILLER_0_23_8 ();
 sg13g2_fill_8 FILLER_0_23_16 ();
 sg13g2_fill_8 FILLER_0_23_24 ();
 sg13g2_fill_2 FILLER_0_23_32 ();
 sg13g2_fill_1 FILLER_0_23_34 ();
 sg13g2_fill_2 FILLER_0_23_61 ();
 sg13g2_fill_1 FILLER_0_23_63 ();
 sg13g2_fill_4 FILLER_0_23_74 ();
 sg13g2_fill_2 FILLER_0_23_78 ();
 sg13g2_fill_2 FILLER_0_23_106 ();
 sg13g2_fill_2 FILLER_0_23_113 ();
 sg13g2_fill_2 FILLER_0_23_120 ();
 sg13g2_fill_2 FILLER_0_23_126 ();
 sg13g2_fill_4 FILLER_0_23_133 ();
 sg13g2_fill_2 FILLER_0_23_137 ();
 sg13g2_fill_2 FILLER_0_23_165 ();
 sg13g2_fill_1 FILLER_0_23_167 ();
 sg13g2_fill_4 FILLER_0_23_178 ();
 sg13g2_fill_4 FILLER_0_23_186 ();
 sg13g2_fill_1 FILLER_0_23_190 ();
 sg13g2_fill_4 FILLER_0_23_195 ();
 sg13g2_fill_1 FILLER_0_23_199 ();
 sg13g2_fill_4 FILLER_0_23_205 ();
 sg13g2_fill_8 FILLER_0_23_213 ();
 sg13g2_fill_8 FILLER_0_23_225 ();
 sg13g2_fill_2 FILLER_0_23_233 ();
 sg13g2_fill_4 FILLER_0_23_239 ();
 sg13g2_fill_4 FILLER_0_23_247 ();
 sg13g2_fill_1 FILLER_0_23_251 ();
 sg13g2_fill_2 FILLER_0_23_258 ();
 sg13g2_fill_2 FILLER_0_23_268 ();
 sg13g2_fill_8 FILLER_0_23_275 ();
 sg13g2_fill_1 FILLER_0_23_283 ();
 sg13g2_fill_4 FILLER_0_23_291 ();
 sg13g2_fill_2 FILLER_0_23_321 ();
 sg13g2_fill_8 FILLER_0_24_0 ();
 sg13g2_fill_8 FILLER_0_24_8 ();
 sg13g2_fill_8 FILLER_0_24_16 ();
 sg13g2_fill_2 FILLER_0_24_34 ();
 sg13g2_fill_4 FILLER_0_24_62 ();
 sg13g2_fill_1 FILLER_0_24_66 ();
 sg13g2_fill_2 FILLER_0_24_93 ();
 sg13g2_fill_4 FILLER_0_24_99 ();
 sg13g2_fill_1 FILLER_0_24_103 ();
 sg13g2_fill_4 FILLER_0_24_109 ();
 sg13g2_fill_2 FILLER_0_24_118 ();
 sg13g2_fill_2 FILLER_0_24_127 ();
 sg13g2_fill_1 FILLER_0_24_129 ();
 sg13g2_fill_4 FILLER_0_24_156 ();
 sg13g2_fill_4 FILLER_0_24_164 ();
 sg13g2_fill_2 FILLER_0_24_168 ();
 sg13g2_fill_4 FILLER_0_24_175 ();
 sg13g2_fill_4 FILLER_0_24_184 ();
 sg13g2_fill_2 FILLER_0_24_188 ();
 sg13g2_fill_4 FILLER_0_24_195 ();
 sg13g2_fill_2 FILLER_0_24_199 ();
 sg13g2_fill_4 FILLER_0_24_227 ();
 sg13g2_fill_1 FILLER_0_24_231 ();
 sg13g2_fill_2 FILLER_0_24_236 ();
 sg13g2_fill_2 FILLER_0_24_243 ();
 sg13g2_fill_8 FILLER_0_24_249 ();
 sg13g2_fill_8 FILLER_0_24_257 ();
 sg13g2_fill_2 FILLER_0_24_271 ();
 sg13g2_fill_1 FILLER_0_24_273 ();
 sg13g2_fill_2 FILLER_0_24_279 ();
 sg13g2_fill_2 FILLER_0_24_286 ();
 sg13g2_fill_1 FILLER_0_24_288 ();
 sg13g2_fill_2 FILLER_0_24_298 ();
 sg13g2_fill_1 FILLER_0_24_300 ();
 sg13g2_fill_4 FILLER_0_24_309 ();
 sg13g2_fill_4 FILLER_0_24_318 ();
 sg13g2_fill_1 FILLER_0_24_322 ();
 sg13g2_fill_8 FILLER_0_25_0 ();
 sg13g2_fill_8 FILLER_0_25_8 ();
 sg13g2_fill_8 FILLER_0_25_16 ();
 sg13g2_fill_8 FILLER_0_25_24 ();
 sg13g2_fill_2 FILLER_0_25_32 ();
 sg13g2_fill_2 FILLER_0_25_38 ();
 sg13g2_fill_2 FILLER_0_25_44 ();
 sg13g2_fill_2 FILLER_0_25_56 ();
 sg13g2_fill_2 FILLER_0_25_84 ();
 sg13g2_fill_2 FILLER_0_25_90 ();
 sg13g2_fill_4 FILLER_0_25_96 ();
 sg13g2_fill_2 FILLER_0_25_100 ();
 sg13g2_fill_4 FILLER_0_25_107 ();
 sg13g2_fill_2 FILLER_0_25_111 ();
 sg13g2_fill_4 FILLER_0_25_118 ();
 sg13g2_fill_4 FILLER_0_25_126 ();
 sg13g2_fill_2 FILLER_0_25_130 ();
 sg13g2_fill_2 FILLER_0_25_158 ();
 sg13g2_fill_1 FILLER_0_25_160 ();
 sg13g2_fill_2 FILLER_0_25_187 ();
 sg13g2_fill_1 FILLER_0_25_189 ();
 sg13g2_fill_2 FILLER_0_25_198 ();
 sg13g2_fill_2 FILLER_0_25_205 ();
 sg13g2_fill_1 FILLER_0_25_207 ();
 sg13g2_fill_2 FILLER_0_25_215 ();
 sg13g2_fill_1 FILLER_0_25_217 ();
 sg13g2_fill_8 FILLER_0_25_222 ();
 sg13g2_fill_2 FILLER_0_25_230 ();
 sg13g2_fill_2 FILLER_0_25_239 ();
 sg13g2_fill_2 FILLER_0_25_246 ();
 sg13g2_fill_2 FILLER_0_25_253 ();
 sg13g2_fill_2 FILLER_0_25_260 ();
 sg13g2_fill_1 FILLER_0_25_262 ();
 sg13g2_fill_2 FILLER_0_25_268 ();
 sg13g2_fill_2 FILLER_0_25_275 ();
 sg13g2_fill_2 FILLER_0_25_281 ();
 sg13g2_fill_2 FILLER_0_25_289 ();
 sg13g2_fill_2 FILLER_0_25_295 ();
 sg13g2_fill_4 FILLER_0_25_307 ();
 sg13g2_fill_2 FILLER_0_25_321 ();
 sg13g2_fill_2 FILLER_0_26_0 ();
 sg13g2_fill_1 FILLER_0_26_2 ();
 sg13g2_fill_4 FILLER_0_26_29 ();
 sg13g2_fill_1 FILLER_0_26_33 ();
 sg13g2_fill_2 FILLER_0_26_38 ();
 sg13g2_fill_1 FILLER_0_26_40 ();
 sg13g2_fill_8 FILLER_0_26_44 ();
 sg13g2_fill_2 FILLER_0_26_52 ();
 sg13g2_fill_1 FILLER_0_26_54 ();
 sg13g2_fill_2 FILLER_0_26_59 ();
 sg13g2_fill_2 FILLER_0_26_87 ();
 sg13g2_fill_8 FILLER_0_26_93 ();
 sg13g2_fill_2 FILLER_0_26_109 ();
 sg13g2_fill_2 FILLER_0_26_115 ();
 sg13g2_fill_1 FILLER_0_26_117 ();
 sg13g2_fill_2 FILLER_0_26_123 ();
 sg13g2_fill_1 FILLER_0_26_125 ();
 sg13g2_fill_4 FILLER_0_26_132 ();
 sg13g2_fill_2 FILLER_0_26_140 ();
 sg13g2_fill_4 FILLER_0_26_168 ();
 sg13g2_fill_4 FILLER_0_26_176 ();
 sg13g2_fill_1 FILLER_0_26_180 ();
 sg13g2_fill_2 FILLER_0_26_186 ();
 sg13g2_fill_2 FILLER_0_26_195 ();
 sg13g2_fill_2 FILLER_0_26_201 ();
 sg13g2_fill_2 FILLER_0_26_229 ();
 sg13g2_fill_2 FILLER_0_26_236 ();
 sg13g2_fill_8 FILLER_0_26_242 ();
 sg13g2_fill_4 FILLER_0_26_250 ();
 sg13g2_fill_1 FILLER_0_26_254 ();
 sg13g2_fill_2 FILLER_0_26_259 ();
 sg13g2_fill_2 FILLER_0_26_266 ();
 sg13g2_fill_2 FILLER_0_26_272 ();
 sg13g2_fill_2 FILLER_0_26_280 ();
 sg13g2_fill_2 FILLER_0_26_287 ();
 sg13g2_fill_8 FILLER_0_26_294 ();
 sg13g2_fill_2 FILLER_0_26_307 ();
 sg13g2_fill_2 FILLER_0_26_314 ();
 sg13g2_fill_2 FILLER_0_26_321 ();
 sg13g2_fill_8 FILLER_0_27_0 ();
 sg13g2_fill_1 FILLER_0_27_8 ();
 sg13g2_fill_8 FILLER_0_27_13 ();
 sg13g2_fill_4 FILLER_0_27_21 ();
 sg13g2_fill_1 FILLER_0_27_25 ();
 sg13g2_fill_4 FILLER_0_27_52 ();
 sg13g2_fill_4 FILLER_0_27_66 ();
 sg13g2_fill_1 FILLER_0_27_70 ();
 sg13g2_fill_8 FILLER_0_27_75 ();
 sg13g2_fill_4 FILLER_0_27_83 ();
 sg13g2_fill_2 FILLER_0_27_87 ();
 sg13g2_fill_2 FILLER_0_27_97 ();
 sg13g2_fill_2 FILLER_0_27_105 ();
 sg13g2_fill_2 FILLER_0_27_115 ();
 sg13g2_fill_2 FILLER_0_27_122 ();
 sg13g2_fill_1 FILLER_0_27_124 ();
 sg13g2_fill_2 FILLER_0_27_128 ();
 sg13g2_fill_2 FILLER_0_27_134 ();
 sg13g2_fill_2 FILLER_0_27_140 ();
 sg13g2_fill_4 FILLER_0_27_168 ();
 sg13g2_fill_8 FILLER_0_27_176 ();
 sg13g2_fill_4 FILLER_0_27_184 ();
 sg13g2_fill_1 FILLER_0_27_188 ();
 sg13g2_fill_2 FILLER_0_27_193 ();
 sg13g2_fill_4 FILLER_0_27_198 ();
 sg13g2_fill_2 FILLER_0_27_228 ();
 sg13g2_fill_2 FILLER_0_27_256 ();
 sg13g2_fill_2 FILLER_0_27_262 ();
 sg13g2_fill_2 FILLER_0_27_268 ();
 sg13g2_fill_1 FILLER_0_27_270 ();
 sg13g2_fill_2 FILLER_0_27_277 ();
 sg13g2_fill_2 FILLER_0_27_283 ();
 sg13g2_fill_1 FILLER_0_27_285 ();
 sg13g2_fill_2 FILLER_0_27_293 ();
 sg13g2_fill_2 FILLER_0_27_300 ();
 sg13g2_fill_2 FILLER_0_27_309 ();
 sg13g2_fill_4 FILLER_0_27_316 ();
 sg13g2_fill_2 FILLER_0_27_320 ();
 sg13g2_fill_1 FILLER_0_27_322 ();
 sg13g2_fill_8 FILLER_0_28_0 ();
 sg13g2_fill_1 FILLER_0_28_8 ();
 sg13g2_fill_2 FILLER_0_28_13 ();
 sg13g2_fill_1 FILLER_0_28_15 ();
 sg13g2_fill_2 FILLER_0_28_24 ();
 sg13g2_fill_2 FILLER_0_28_30 ();
 sg13g2_fill_2 FILLER_0_28_40 ();
 sg13g2_fill_2 FILLER_0_28_46 ();
 sg13g2_fill_8 FILLER_0_28_52 ();
 sg13g2_fill_4 FILLER_0_28_60 ();
 sg13g2_fill_2 FILLER_0_28_64 ();
 sg13g2_fill_1 FILLER_0_28_66 ();
 sg13g2_fill_2 FILLER_0_28_93 ();
 sg13g2_fill_4 FILLER_0_28_100 ();
 sg13g2_fill_4 FILLER_0_28_111 ();
 sg13g2_fill_2 FILLER_0_28_115 ();
 sg13g2_fill_2 FILLER_0_28_122 ();
 sg13g2_fill_2 FILLER_0_28_129 ();
 sg13g2_fill_2 FILLER_0_28_135 ();
 sg13g2_fill_4 FILLER_0_28_142 ();
 sg13g2_fill_2 FILLER_0_28_146 ();
 sg13g2_fill_2 FILLER_0_28_152 ();
 sg13g2_fill_2 FILLER_0_28_158 ();
 sg13g2_fill_2 FILLER_0_28_164 ();
 sg13g2_fill_2 FILLER_0_28_192 ();
 sg13g2_fill_4 FILLER_0_28_199 ();
 sg13g2_fill_2 FILLER_0_28_207 ();
 sg13g2_fill_4 FILLER_0_28_213 ();
 sg13g2_fill_4 FILLER_0_28_221 ();
 sg13g2_fill_4 FILLER_0_28_230 ();
 sg13g2_fill_2 FILLER_0_28_234 ();
 sg13g2_fill_4 FILLER_0_28_240 ();
 sg13g2_fill_2 FILLER_0_28_244 ();
 sg13g2_fill_4 FILLER_0_28_250 ();
 sg13g2_fill_2 FILLER_0_28_254 ();
 sg13g2_fill_2 FILLER_0_28_261 ();
 sg13g2_fill_1 FILLER_0_28_263 ();
 sg13g2_fill_2 FILLER_0_28_272 ();
 sg13g2_fill_2 FILLER_0_28_277 ();
 sg13g2_fill_2 FILLER_0_28_286 ();
 sg13g2_fill_2 FILLER_0_28_296 ();
 sg13g2_fill_2 FILLER_0_28_305 ();
 sg13g2_fill_2 FILLER_0_28_314 ();
 sg13g2_fill_1 FILLER_0_28_316 ();
 sg13g2_fill_1 FILLER_0_28_322 ();
 sg13g2_fill_4 FILLER_0_29_0 ();
 sg13g2_fill_2 FILLER_0_29_4 ();
 sg13g2_fill_1 FILLER_0_29_6 ();
 sg13g2_fill_2 FILLER_0_29_11 ();
 sg13g2_fill_1 FILLER_0_29_13 ();
 sg13g2_fill_2 FILLER_0_29_18 ();
 sg13g2_fill_2 FILLER_0_29_28 ();
 sg13g2_fill_4 FILLER_0_29_34 ();
 sg13g2_fill_2 FILLER_0_29_46 ();
 sg13g2_fill_2 FILLER_0_29_74 ();
 sg13g2_fill_1 FILLER_0_29_76 ();
 sg13g2_fill_4 FILLER_0_29_81 ();
 sg13g2_fill_4 FILLER_0_29_89 ();
 sg13g2_fill_4 FILLER_0_29_97 ();
 sg13g2_fill_2 FILLER_0_29_106 ();
 sg13g2_fill_8 FILLER_0_29_116 ();
 sg13g2_fill_8 FILLER_0_29_124 ();
 sg13g2_fill_2 FILLER_0_29_132 ();
 sg13g2_fill_1 FILLER_0_29_134 ();
 sg13g2_fill_8 FILLER_0_29_161 ();
 sg13g2_fill_2 FILLER_0_29_169 ();
 sg13g2_fill_8 FILLER_0_29_175 ();
 sg13g2_fill_8 FILLER_0_29_183 ();
 sg13g2_fill_2 FILLER_0_29_196 ();
 sg13g2_fill_2 FILLER_0_29_205 ();
 sg13g2_fill_1 FILLER_0_29_207 ();
 sg13g2_fill_4 FILLER_0_29_234 ();
 sg13g2_fill_2 FILLER_0_29_238 ();
 sg13g2_fill_2 FILLER_0_29_245 ();
 sg13g2_fill_1 FILLER_0_29_247 ();
 sg13g2_fill_2 FILLER_0_29_256 ();
 sg13g2_fill_1 FILLER_0_29_258 ();
 sg13g2_fill_2 FILLER_0_29_263 ();
 sg13g2_fill_1 FILLER_0_29_265 ();
 sg13g2_fill_4 FILLER_0_29_274 ();
 sg13g2_fill_2 FILLER_0_29_283 ();
 sg13g2_fill_2 FILLER_0_29_290 ();
 sg13g2_fill_8 FILLER_0_29_298 ();
 sg13g2_fill_4 FILLER_0_29_316 ();
 sg13g2_fill_2 FILLER_0_29_320 ();
 sg13g2_fill_1 FILLER_0_29_322 ();
 sg13g2_fill_4 FILLER_0_30_0 ();
 sg13g2_fill_1 FILLER_0_30_4 ();
 sg13g2_fill_2 FILLER_0_30_31 ();
 sg13g2_fill_4 FILLER_0_30_38 ();
 sg13g2_fill_2 FILLER_0_30_42 ();
 sg13g2_fill_1 FILLER_0_30_44 ();
 sg13g2_fill_4 FILLER_0_30_50 ();
 sg13g2_fill_2 FILLER_0_30_54 ();
 sg13g2_fill_4 FILLER_0_30_60 ();
 sg13g2_fill_2 FILLER_0_30_64 ();
 sg13g2_fill_4 FILLER_0_30_92 ();
 sg13g2_fill_2 FILLER_0_30_96 ();
 sg13g2_fill_2 FILLER_0_30_106 ();
 sg13g2_fill_4 FILLER_0_30_113 ();
 sg13g2_fill_1 FILLER_0_30_117 ();
 sg13g2_fill_2 FILLER_0_30_125 ();
 sg13g2_fill_4 FILLER_0_30_133 ();
 sg13g2_fill_1 FILLER_0_30_137 ();
 sg13g2_fill_2 FILLER_0_30_164 ();
 sg13g2_fill_2 FILLER_0_30_192 ();
 sg13g2_fill_2 FILLER_0_30_198 ();
 sg13g2_fill_2 FILLER_0_30_210 ();
 sg13g2_fill_2 FILLER_0_30_217 ();
 sg13g2_fill_4 FILLER_0_30_224 ();
 sg13g2_fill_4 FILLER_0_30_254 ();
 sg13g2_fill_1 FILLER_0_30_258 ();
 sg13g2_fill_4 FILLER_0_30_265 ();
 sg13g2_fill_1 FILLER_0_30_269 ();
 sg13g2_fill_4 FILLER_0_30_278 ();
 sg13g2_fill_1 FILLER_0_30_282 ();
 sg13g2_fill_8 FILLER_0_30_291 ();
 sg13g2_fill_4 FILLER_0_30_299 ();
 sg13g2_fill_2 FILLER_0_30_309 ();
 sg13g2_fill_4 FILLER_0_30_317 ();
 sg13g2_fill_2 FILLER_0_30_321 ();
 sg13g2_fill_2 FILLER_0_31_0 ();
 sg13g2_fill_1 FILLER_0_31_2 ();
 sg13g2_fill_2 FILLER_0_31_29 ();
 sg13g2_fill_4 FILLER_0_31_37 ();
 sg13g2_fill_1 FILLER_0_31_41 ();
 sg13g2_fill_2 FILLER_0_31_50 ();
 sg13g2_fill_2 FILLER_0_31_78 ();
 sg13g2_fill_1 FILLER_0_31_80 ();
 sg13g2_fill_2 FILLER_0_31_89 ();
 sg13g2_fill_2 FILLER_0_31_96 ();
 sg13g2_fill_2 FILLER_0_31_106 ();
 sg13g2_fill_1 FILLER_0_31_108 ();
 sg13g2_fill_2 FILLER_0_31_114 ();
 sg13g2_fill_1 FILLER_0_31_116 ();
 sg13g2_fill_2 FILLER_0_31_120 ();
 sg13g2_fill_2 FILLER_0_31_127 ();
 sg13g2_fill_2 FILLER_0_31_132 ();
 sg13g2_fill_2 FILLER_0_31_140 ();
 sg13g2_fill_2 FILLER_0_31_146 ();
 sg13g2_fill_2 FILLER_0_31_152 ();
 sg13g2_fill_4 FILLER_0_31_158 ();
 sg13g2_fill_4 FILLER_0_31_167 ();
 sg13g2_fill_2 FILLER_0_31_174 ();
 sg13g2_fill_1 FILLER_0_31_176 ();
 sg13g2_fill_2 FILLER_0_31_181 ();
 sg13g2_fill_1 FILLER_0_31_183 ();
 sg13g2_fill_4 FILLER_0_31_189 ();
 sg13g2_fill_2 FILLER_0_31_198 ();
 sg13g2_fill_4 FILLER_0_31_204 ();
 sg13g2_fill_2 FILLER_0_31_208 ();
 sg13g2_fill_4 FILLER_0_31_215 ();
 sg13g2_fill_2 FILLER_0_31_224 ();
 sg13g2_fill_1 FILLER_0_31_226 ();
 sg13g2_fill_4 FILLER_0_31_232 ();
 sg13g2_fill_2 FILLER_0_31_236 ();
 sg13g2_fill_1 FILLER_0_31_238 ();
 sg13g2_fill_8 FILLER_0_31_244 ();
 sg13g2_fill_4 FILLER_0_31_252 ();
 sg13g2_fill_2 FILLER_0_31_256 ();
 sg13g2_fill_4 FILLER_0_31_266 ();
 sg13g2_fill_1 FILLER_0_31_270 ();
 sg13g2_fill_2 FILLER_0_31_277 ();
 sg13g2_fill_4 FILLER_0_31_288 ();
 sg13g2_fill_2 FILLER_0_31_292 ();
 sg13g2_fill_1 FILLER_0_31_294 ();
 sg13g2_fill_2 FILLER_0_31_321 ();
 sg13g2_fill_1 FILLER_0_32_0 ();
 sg13g2_fill_2 FILLER_0_32_5 ();
 sg13g2_fill_2 FILLER_0_32_11 ();
 sg13g2_fill_2 FILLER_0_32_21 ();
 sg13g2_fill_2 FILLER_0_32_27 ();
 sg13g2_fill_8 FILLER_0_32_32 ();
 sg13g2_fill_2 FILLER_0_32_46 ();
 sg13g2_fill_2 FILLER_0_32_52 ();
 sg13g2_fill_4 FILLER_0_32_62 ();
 sg13g2_fill_2 FILLER_0_32_66 ();
 sg13g2_fill_4 FILLER_0_32_72 ();
 sg13g2_fill_4 FILLER_0_32_80 ();
 sg13g2_fill_4 FILLER_0_32_88 ();
 sg13g2_fill_4 FILLER_0_32_97 ();
 sg13g2_fill_4 FILLER_0_32_104 ();
 sg13g2_fill_1 FILLER_0_32_108 ();
 sg13g2_fill_8 FILLER_0_32_114 ();
 sg13g2_fill_4 FILLER_0_32_122 ();
 sg13g2_fill_2 FILLER_0_32_126 ();
 sg13g2_fill_1 FILLER_0_32_128 ();
 sg13g2_fill_2 FILLER_0_32_134 ();
 sg13g2_fill_4 FILLER_0_32_141 ();
 sg13g2_fill_2 FILLER_0_32_145 ();
 sg13g2_fill_1 FILLER_0_32_147 ();
 sg13g2_fill_2 FILLER_0_32_152 ();
 sg13g2_fill_2 FILLER_0_32_159 ();
 sg13g2_fill_1 FILLER_0_32_161 ();
 sg13g2_fill_2 FILLER_0_32_168 ();
 sg13g2_fill_4 FILLER_0_32_176 ();
 sg13g2_fill_4 FILLER_0_32_185 ();
 sg13g2_fill_1 FILLER_0_32_189 ();
 sg13g2_fill_4 FILLER_0_32_193 ();
 sg13g2_fill_2 FILLER_0_32_197 ();
 sg13g2_fill_4 FILLER_0_32_204 ();
 sg13g2_fill_4 FILLER_0_32_211 ();
 sg13g2_fill_2 FILLER_0_32_215 ();
 sg13g2_fill_1 FILLER_0_32_217 ();
 sg13g2_fill_2 FILLER_0_32_223 ();
 sg13g2_fill_4 FILLER_0_32_251 ();
 sg13g2_fill_2 FILLER_0_32_255 ();
 sg13g2_fill_2 FILLER_0_32_262 ();
 sg13g2_fill_2 FILLER_0_32_269 ();
 sg13g2_fill_2 FILLER_0_32_276 ();
 sg13g2_fill_2 FILLER_0_32_283 ();
 sg13g2_fill_8 FILLER_0_32_290 ();
 sg13g2_fill_2 FILLER_0_32_302 ();
 sg13g2_fill_4 FILLER_0_32_308 ();
 sg13g2_fill_2 FILLER_0_32_320 ();
 sg13g2_fill_1 FILLER_0_32_322 ();
 sg13g2_fill_4 FILLER_0_33_0 ();
 sg13g2_fill_2 FILLER_0_33_4 ();
 sg13g2_fill_1 FILLER_0_33_6 ();
 sg13g2_fill_4 FILLER_0_33_11 ();
 sg13g2_fill_4 FILLER_0_33_23 ();
 sg13g2_fill_2 FILLER_0_33_30 ();
 sg13g2_fill_2 FILLER_0_33_41 ();
 sg13g2_fill_1 FILLER_0_33_43 ();
 sg13g2_fill_2 FILLER_0_33_48 ();
 sg13g2_fill_4 FILLER_0_33_76 ();
 sg13g2_fill_2 FILLER_0_33_80 ();
 sg13g2_fill_2 FILLER_0_33_90 ();
 sg13g2_fill_4 FILLER_0_33_97 ();
 sg13g2_fill_2 FILLER_0_33_101 ();
 sg13g2_fill_4 FILLER_0_33_107 ();
 sg13g2_fill_4 FILLER_0_33_116 ();
 sg13g2_fill_1 FILLER_0_33_120 ();
 sg13g2_fill_4 FILLER_0_33_127 ();
 sg13g2_fill_4 FILLER_0_33_136 ();
 sg13g2_fill_2 FILLER_0_33_140 ();
 sg13g2_fill_4 FILLER_0_33_147 ();
 sg13g2_fill_2 FILLER_0_33_177 ();
 sg13g2_fill_4 FILLER_0_33_184 ();
 sg13g2_fill_2 FILLER_0_33_191 ();
 sg13g2_fill_2 FILLER_0_33_203 ();
 sg13g2_fill_2 FILLER_0_33_231 ();
 sg13g2_fill_2 FILLER_0_33_237 ();
 sg13g2_fill_2 FILLER_0_33_265 ();
 sg13g2_fill_2 FILLER_0_33_272 ();
 sg13g2_fill_2 FILLER_0_33_279 ();
 sg13g2_fill_1 FILLER_0_33_281 ();
 sg13g2_fill_2 FILLER_0_33_287 ();
 sg13g2_fill_2 FILLER_0_33_293 ();
 sg13g2_fill_2 FILLER_0_33_321 ();
 sg13g2_fill_4 FILLER_0_34_0 ();
 sg13g2_fill_4 FILLER_0_34_30 ();
 sg13g2_fill_1 FILLER_0_34_34 ();
 sg13g2_fill_2 FILLER_0_34_43 ();
 sg13g2_fill_1 FILLER_0_34_45 ();
 sg13g2_fill_2 FILLER_0_34_50 ();
 sg13g2_fill_1 FILLER_0_34_52 ();
 sg13g2_fill_4 FILLER_0_34_58 ();
 sg13g2_fill_4 FILLER_0_34_66 ();
 sg13g2_fill_2 FILLER_0_34_96 ();
 sg13g2_fill_1 FILLER_0_34_98 ();
 sg13g2_fill_2 FILLER_0_34_103 ();
 sg13g2_fill_1 FILLER_0_34_105 ();
 sg13g2_fill_4 FILLER_0_34_111 ();
 sg13g2_fill_2 FILLER_0_34_120 ();
 sg13g2_fill_1 FILLER_0_34_122 ();
 sg13g2_fill_4 FILLER_0_34_131 ();
 sg13g2_fill_2 FILLER_0_34_140 ();
 sg13g2_fill_1 FILLER_0_34_142 ();
 sg13g2_fill_2 FILLER_0_34_148 ();
 sg13g2_fill_1 FILLER_0_34_150 ();
 sg13g2_fill_2 FILLER_0_34_156 ();
 sg13g2_fill_1 FILLER_0_34_158 ();
 sg13g2_fill_2 FILLER_0_34_163 ();
 sg13g2_fill_1 FILLER_0_34_165 ();
 sg13g2_fill_2 FILLER_0_34_171 ();
 sg13g2_fill_1 FILLER_0_34_173 ();
 sg13g2_fill_2 FILLER_0_34_179 ();
 sg13g2_fill_2 FILLER_0_34_185 ();
 sg13g2_fill_2 FILLER_0_34_191 ();
 sg13g2_fill_4 FILLER_0_34_197 ();
 sg13g2_fill_4 FILLER_0_34_206 ();
 sg13g2_fill_2 FILLER_0_34_210 ();
 sg13g2_fill_2 FILLER_0_34_216 ();
 sg13g2_fill_1 FILLER_0_34_218 ();
 sg13g2_fill_2 FILLER_0_34_224 ();
 sg13g2_fill_1 FILLER_0_34_226 ();
 sg13g2_fill_2 FILLER_0_34_253 ();
 sg13g2_fill_2 FILLER_0_34_260 ();
 sg13g2_fill_4 FILLER_0_34_267 ();
 sg13g2_fill_2 FILLER_0_34_271 ();
 sg13g2_fill_1 FILLER_0_34_273 ();
 sg13g2_fill_2 FILLER_0_34_282 ();
 sg13g2_fill_1 FILLER_0_34_284 ();
 sg13g2_fill_2 FILLER_0_34_290 ();
 sg13g2_fill_2 FILLER_0_34_297 ();
 sg13g2_fill_8 FILLER_0_34_303 ();
 sg13g2_fill_2 FILLER_0_34_311 ();
 sg13g2_fill_4 FILLER_0_34_317 ();
 sg13g2_fill_2 FILLER_0_34_321 ();
 sg13g2_fill_2 FILLER_0_35_0 ();
 sg13g2_fill_1 FILLER_0_35_2 ();
 sg13g2_fill_4 FILLER_0_35_7 ();
 sg13g2_fill_1 FILLER_0_35_11 ();
 sg13g2_fill_4 FILLER_0_35_16 ();
 sg13g2_fill_1 FILLER_0_35_20 ();
 sg13g2_fill_4 FILLER_0_35_25 ();
 sg13g2_fill_4 FILLER_0_35_34 ();
 sg13g2_fill_1 FILLER_0_35_38 ();
 sg13g2_fill_2 FILLER_0_35_43 ();
 sg13g2_fill_4 FILLER_0_35_71 ();
 sg13g2_fill_2 FILLER_0_35_101 ();
 sg13g2_fill_2 FILLER_0_35_109 ();
 sg13g2_fill_2 FILLER_0_35_116 ();
 sg13g2_fill_2 FILLER_0_35_124 ();
 sg13g2_fill_2 FILLER_0_35_131 ();
 sg13g2_fill_4 FILLER_0_35_136 ();
 sg13g2_fill_2 FILLER_0_35_140 ();
 sg13g2_fill_1 FILLER_0_35_142 ();
 sg13g2_fill_2 FILLER_0_35_148 ();
 sg13g2_fill_2 FILLER_0_35_155 ();
 sg13g2_fill_2 FILLER_0_35_160 ();
 sg13g2_fill_2 FILLER_0_35_188 ();
 sg13g2_fill_2 FILLER_0_35_198 ();
 sg13g2_fill_2 FILLER_0_35_204 ();
 sg13g2_fill_2 FILLER_0_35_210 ();
 sg13g2_fill_2 FILLER_0_35_216 ();
 sg13g2_fill_2 FILLER_0_35_226 ();
 sg13g2_fill_1 FILLER_0_35_228 ();
 sg13g2_fill_2 FILLER_0_35_234 ();
 sg13g2_fill_2 FILLER_0_35_240 ();
 sg13g2_fill_1 FILLER_0_35_242 ();
 sg13g2_fill_2 FILLER_0_35_247 ();
 sg13g2_fill_1 FILLER_0_35_249 ();
 sg13g2_fill_2 FILLER_0_35_255 ();
 sg13g2_fill_2 FILLER_0_35_261 ();
 sg13g2_fill_4 FILLER_0_35_267 ();
 sg13g2_fill_1 FILLER_0_35_271 ();
 sg13g2_fill_2 FILLER_0_35_277 ();
 sg13g2_fill_8 FILLER_0_35_286 ();
 sg13g2_fill_2 FILLER_0_35_294 ();
 sg13g2_fill_4 FILLER_0_35_300 ();
 sg13g2_fill_4 FILLER_0_35_308 ();
 sg13g2_fill_4 FILLER_0_35_317 ();
 sg13g2_fill_2 FILLER_0_35_321 ();
 sg13g2_fill_1 FILLER_0_36_0 ();
 sg13g2_fill_2 FILLER_0_36_5 ();
 sg13g2_fill_2 FILLER_0_36_33 ();
 sg13g2_fill_4 FILLER_0_36_40 ();
 sg13g2_fill_2 FILLER_0_36_48 ();
 sg13g2_fill_4 FILLER_0_36_76 ();
 sg13g2_fill_2 FILLER_0_36_84 ();
 sg13g2_fill_2 FILLER_0_36_96 ();
 sg13g2_fill_1 FILLER_0_36_98 ();
 sg13g2_fill_2 FILLER_0_36_103 ();
 sg13g2_fill_1 FILLER_0_36_105 ();
 sg13g2_fill_4 FILLER_0_36_111 ();
 sg13g2_fill_1 FILLER_0_36_115 ();
 sg13g2_fill_2 FILLER_0_36_121 ();
 sg13g2_fill_2 FILLER_0_36_127 ();
 sg13g2_fill_4 FILLER_0_36_134 ();
 sg13g2_fill_2 FILLER_0_36_143 ();
 sg13g2_fill_1 FILLER_0_36_145 ();
 sg13g2_fill_2 FILLER_0_36_150 ();
 sg13g2_fill_1 FILLER_0_36_152 ();
 sg13g2_fill_2 FILLER_0_36_160 ();
 sg13g2_fill_1 FILLER_0_36_162 ();
 sg13g2_fill_2 FILLER_0_36_168 ();
 sg13g2_fill_1 FILLER_0_36_170 ();
 sg13g2_fill_2 FILLER_0_36_175 ();
 sg13g2_fill_1 FILLER_0_36_177 ();
 sg13g2_fill_2 FILLER_0_36_183 ();
 sg13g2_fill_1 FILLER_0_36_185 ();
 sg13g2_fill_2 FILLER_0_36_191 ();
 sg13g2_fill_2 FILLER_0_36_202 ();
 sg13g2_fill_2 FILLER_0_36_209 ();
 sg13g2_fill_2 FILLER_0_36_215 ();
 sg13g2_fill_1 FILLER_0_36_217 ();
 sg13g2_fill_4 FILLER_0_36_222 ();
 sg13g2_fill_2 FILLER_0_36_231 ();
 sg13g2_fill_2 FILLER_0_36_238 ();
 sg13g2_fill_2 FILLER_0_36_245 ();
 sg13g2_fill_4 FILLER_0_36_252 ();
 sg13g2_fill_2 FILLER_0_36_256 ();
 sg13g2_fill_1 FILLER_0_36_258 ();
 sg13g2_fill_2 FILLER_0_36_265 ();
 sg13g2_fill_2 FILLER_0_36_271 ();
 sg13g2_fill_8 FILLER_0_36_278 ();
 sg13g2_fill_2 FILLER_0_36_286 ();
 sg13g2_fill_1 FILLER_0_36_288 ();
 sg13g2_fill_2 FILLER_0_36_293 ();
 sg13g2_fill_2 FILLER_0_36_321 ();
 sg13g2_fill_2 FILLER_0_37_0 ();
 sg13g2_fill_2 FILLER_0_37_10 ();
 sg13g2_fill_1 FILLER_0_37_12 ();
 sg13g2_fill_2 FILLER_0_37_17 ();
 sg13g2_fill_1 FILLER_0_37_19 ();
 sg13g2_fill_4 FILLER_0_37_27 ();
 sg13g2_fill_2 FILLER_0_37_37 ();
 sg13g2_fill_2 FILLER_0_37_45 ();
 sg13g2_fill_2 FILLER_0_37_51 ();
 sg13g2_fill_4 FILLER_0_37_61 ();
 sg13g2_fill_2 FILLER_0_37_69 ();
 sg13g2_fill_4 FILLER_0_37_97 ();
 sg13g2_fill_2 FILLER_0_37_105 ();
 sg13g2_fill_4 FILLER_0_37_112 ();
 sg13g2_fill_2 FILLER_0_37_116 ();
 sg13g2_fill_2 FILLER_0_37_122 ();
 sg13g2_fill_1 FILLER_0_37_124 ();
 sg13g2_fill_4 FILLER_0_37_128 ();
 sg13g2_fill_1 FILLER_0_37_132 ();
 sg13g2_fill_2 FILLER_0_37_139 ();
 sg13g2_fill_4 FILLER_0_37_167 ();
 sg13g2_fill_1 FILLER_0_37_171 ();
 sg13g2_fill_2 FILLER_0_37_177 ();
 sg13g2_fill_4 FILLER_0_37_184 ();
 sg13g2_fill_2 FILLER_0_37_188 ();
 sg13g2_fill_1 FILLER_0_37_190 ();
 sg13g2_fill_2 FILLER_0_37_201 ();
 sg13g2_fill_2 FILLER_0_37_208 ();
 sg13g2_fill_2 FILLER_0_37_215 ();
 sg13g2_fill_4 FILLER_0_37_223 ();
 sg13g2_fill_1 FILLER_0_37_227 ();
 sg13g2_fill_4 FILLER_0_37_238 ();
 sg13g2_fill_1 FILLER_0_37_242 ();
 sg13g2_fill_2 FILLER_0_37_269 ();
 sg13g2_fill_2 FILLER_0_37_275 ();
 sg13g2_fill_4 FILLER_0_37_282 ();
 sg13g2_fill_2 FILLER_0_37_286 ();
 sg13g2_fill_2 FILLER_0_37_293 ();
 sg13g2_fill_2 FILLER_0_37_300 ();
 sg13g2_fill_2 FILLER_0_37_307 ();
 sg13g2_fill_4 FILLER_0_37_317 ();
 sg13g2_fill_2 FILLER_0_37_321 ();
 sg13g2_fill_2 FILLER_0_38_0 ();
 sg13g2_fill_1 FILLER_0_38_2 ();
 sg13g2_fill_2 FILLER_0_38_29 ();
 sg13g2_fill_2 FILLER_0_38_39 ();
 sg13g2_fill_2 FILLER_0_38_67 ();
 sg13g2_fill_2 FILLER_0_38_73 ();
 sg13g2_fill_2 FILLER_0_38_83 ();
 sg13g2_fill_1 FILLER_0_38_85 ();
 sg13g2_fill_2 FILLER_0_38_91 ();
 sg13g2_fill_2 FILLER_0_38_98 ();
 sg13g2_fill_2 FILLER_0_38_105 ();
 sg13g2_fill_1 FILLER_0_38_107 ();
 sg13g2_fill_2 FILLER_0_38_113 ();
 sg13g2_fill_2 FILLER_0_38_120 ();
 sg13g2_fill_1 FILLER_0_38_122 ();
 sg13g2_fill_2 FILLER_0_38_131 ();
 sg13g2_fill_2 FILLER_0_38_138 ();
 sg13g2_fill_2 FILLER_0_38_145 ();
 sg13g2_fill_1 FILLER_0_38_147 ();
 sg13g2_fill_4 FILLER_0_38_152 ();
 sg13g2_fill_1 FILLER_0_38_156 ();
 sg13g2_fill_4 FILLER_0_38_162 ();
 sg13g2_fill_2 FILLER_0_38_166 ();
 sg13g2_fill_1 FILLER_0_38_168 ();
 sg13g2_fill_2 FILLER_0_38_175 ();
 sg13g2_fill_2 FILLER_0_38_182 ();
 sg13g2_fill_1 FILLER_0_38_184 ();
 sg13g2_fill_4 FILLER_0_38_190 ();
 sg13g2_fill_1 FILLER_0_38_194 ();
 sg13g2_fill_2 FILLER_0_38_201 ();
 sg13g2_fill_2 FILLER_0_38_208 ();
 sg13g2_fill_2 FILLER_0_38_215 ();
 sg13g2_fill_1 FILLER_0_38_217 ();
 sg13g2_fill_2 FILLER_0_38_223 ();
 sg13g2_fill_2 FILLER_0_38_230 ();
 sg13g2_fill_1 FILLER_0_38_232 ();
 sg13g2_fill_2 FILLER_0_38_259 ();
 sg13g2_fill_1 FILLER_0_38_261 ();
 sg13g2_fill_4 FILLER_0_38_267 ();
 sg13g2_fill_2 FILLER_0_38_276 ();
 sg13g2_fill_2 FILLER_0_38_285 ();
 sg13g2_fill_1 FILLER_0_38_287 ();
 sg13g2_fill_2 FILLER_0_38_294 ();
 sg13g2_fill_1 FILLER_0_38_296 ();
 sg13g2_fill_2 FILLER_0_38_305 ();
 sg13g2_fill_2 FILLER_0_38_315 ();
 sg13g2_fill_1 FILLER_0_38_317 ();
 sg13g2_fill_1 FILLER_0_38_322 ();
 sg13g2_fill_4 FILLER_0_39_0 ();
 sg13g2_fill_2 FILLER_0_39_4 ();
 sg13g2_fill_2 FILLER_0_39_10 ();
 sg13g2_fill_2 FILLER_0_39_16 ();
 sg13g2_fill_4 FILLER_0_39_26 ();
 sg13g2_fill_2 FILLER_0_39_34 ();
 sg13g2_fill_2 FILLER_0_39_40 ();
 sg13g2_fill_2 FILLER_0_39_46 ();
 sg13g2_fill_2 FILLER_0_39_52 ();
 sg13g2_fill_2 FILLER_0_39_59 ();
 sg13g2_fill_2 FILLER_0_39_67 ();
 sg13g2_fill_2 FILLER_0_39_74 ();
 sg13g2_fill_2 FILLER_0_39_102 ();
 sg13g2_fill_2 FILLER_0_39_109 ();
 sg13g2_fill_2 FILLER_0_39_116 ();
 sg13g2_fill_2 FILLER_0_39_123 ();
 sg13g2_fill_2 FILLER_0_39_130 ();
 sg13g2_fill_1 FILLER_0_39_132 ();
 sg13g2_fill_2 FILLER_0_39_138 ();
 sg13g2_fill_1 FILLER_0_39_140 ();
 sg13g2_fill_2 FILLER_0_39_148 ();
 sg13g2_fill_4 FILLER_0_39_155 ();
 sg13g2_fill_8 FILLER_0_39_169 ();
 sg13g2_fill_2 FILLER_0_39_177 ();
 sg13g2_fill_1 FILLER_0_39_179 ();
 sg13g2_fill_2 FILLER_0_39_185 ();
 sg13g2_fill_2 FILLER_0_39_191 ();
 sg13g2_fill_2 FILLER_0_39_198 ();
 sg13g2_fill_2 FILLER_0_39_206 ();
 sg13g2_fill_4 FILLER_0_39_213 ();
 sg13g2_fill_2 FILLER_0_39_222 ();
 sg13g2_fill_1 FILLER_0_39_224 ();
 sg13g2_fill_2 FILLER_0_39_230 ();
 sg13g2_fill_1 FILLER_0_39_232 ();
 sg13g2_fill_2 FILLER_0_39_238 ();
 sg13g2_fill_1 FILLER_0_39_240 ();
 sg13g2_fill_2 FILLER_0_39_247 ();
 sg13g2_fill_1 FILLER_0_39_249 ();
 sg13g2_fill_4 FILLER_0_39_254 ();
 sg13g2_fill_4 FILLER_0_39_262 ();
 sg13g2_fill_4 FILLER_0_39_274 ();
 sg13g2_fill_2 FILLER_0_39_283 ();
 sg13g2_fill_2 FILLER_0_39_290 ();
 sg13g2_fill_2 FILLER_0_39_297 ();
 sg13g2_fill_4 FILLER_0_39_304 ();
 sg13g2_fill_8 FILLER_0_39_315 ();
 sg13g2_fill_2 FILLER_0_40_0 ();
 sg13g2_fill_2 FILLER_0_40_28 ();
 sg13g2_fill_2 FILLER_0_40_34 ();
 sg13g2_fill_2 FILLER_0_40_44 ();
 sg13g2_fill_2 FILLER_0_40_49 ();
 sg13g2_fill_2 FILLER_0_40_55 ();
 sg13g2_fill_4 FILLER_0_40_64 ();
 sg13g2_fill_1 FILLER_0_40_68 ();
 sg13g2_fill_2 FILLER_0_40_73 ();
 sg13g2_fill_2 FILLER_0_40_78 ();
 sg13g2_fill_2 FILLER_0_40_84 ();
 sg13g2_fill_4 FILLER_0_40_92 ();
 sg13g2_fill_1 FILLER_0_40_96 ();
 sg13g2_fill_2 FILLER_0_40_102 ();
 sg13g2_fill_2 FILLER_0_40_112 ();
 sg13g2_fill_2 FILLER_0_40_117 ();
 sg13g2_fill_1 FILLER_0_40_119 ();
 sg13g2_fill_2 FILLER_0_40_125 ();
 sg13g2_fill_1 FILLER_0_40_127 ();
 sg13g2_fill_2 FILLER_0_40_133 ();
 sg13g2_fill_2 FILLER_0_40_140 ();
 sg13g2_fill_1 FILLER_0_40_142 ();
 sg13g2_fill_4 FILLER_0_40_169 ();
 sg13g2_fill_4 FILLER_0_40_177 ();
 sg13g2_fill_2 FILLER_0_40_189 ();
 sg13g2_fill_1 FILLER_0_40_191 ();
 sg13g2_fill_2 FILLER_0_40_197 ();
 sg13g2_fill_4 FILLER_0_40_204 ();
 sg13g2_fill_4 FILLER_0_40_213 ();
 sg13g2_fill_2 FILLER_0_40_222 ();
 sg13g2_fill_2 FILLER_0_40_229 ();
 sg13g2_fill_2 FILLER_0_40_235 ();
 sg13g2_fill_2 FILLER_0_40_240 ();
 sg13g2_fill_2 FILLER_0_40_268 ();
 sg13g2_fill_1 FILLER_0_40_270 ();
 sg13g2_fill_4 FILLER_0_40_275 ();
 sg13g2_fill_2 FILLER_0_40_279 ();
 sg13g2_fill_1 FILLER_0_40_281 ();
 sg13g2_fill_2 FILLER_0_40_287 ();
 sg13g2_fill_1 FILLER_0_40_289 ();
 sg13g2_fill_2 FILLER_0_40_296 ();
 sg13g2_fill_4 FILLER_0_40_301 ();
 sg13g2_fill_1 FILLER_0_40_305 ();
 sg13g2_fill_2 FILLER_0_40_313 ();
 sg13g2_fill_4 FILLER_0_40_319 ();
 sg13g2_fill_4 FILLER_0_41_0 ();
 sg13g2_fill_2 FILLER_0_41_30 ();
 sg13g2_fill_2 FILLER_0_41_36 ();
 sg13g2_fill_4 FILLER_0_41_64 ();
 sg13g2_fill_2 FILLER_0_41_68 ();
 sg13g2_fill_1 FILLER_0_41_70 ();
 sg13g2_fill_2 FILLER_0_41_75 ();
 sg13g2_fill_2 FILLER_0_41_83 ();
 sg13g2_fill_2 FILLER_0_41_90 ();
 sg13g2_fill_4 FILLER_0_41_96 ();
 sg13g2_fill_2 FILLER_0_41_104 ();
 sg13g2_fill_1 FILLER_0_41_106 ();
 sg13g2_fill_2 FILLER_0_41_133 ();
 sg13g2_fill_1 FILLER_0_41_135 ();
 sg13g2_fill_2 FILLER_0_41_143 ();
 sg13g2_fill_1 FILLER_0_41_145 ();
 sg13g2_fill_2 FILLER_0_41_150 ();
 sg13g2_fill_1 FILLER_0_41_152 ();
 sg13g2_fill_4 FILLER_0_41_157 ();
 sg13g2_fill_4 FILLER_0_41_165 ();
 sg13g2_fill_4 FILLER_0_41_177 ();
 sg13g2_fill_4 FILLER_0_41_193 ();
 sg13g2_fill_4 FILLER_0_41_202 ();
 sg13g2_fill_2 FILLER_0_41_206 ();
 sg13g2_fill_1 FILLER_0_41_208 ();
 sg13g2_fill_2 FILLER_0_41_215 ();
 sg13g2_fill_2 FILLER_0_41_221 ();
 sg13g2_fill_1 FILLER_0_41_223 ();
 sg13g2_fill_2 FILLER_0_41_231 ();
 sg13g2_fill_2 FILLER_0_41_237 ();
 sg13g2_fill_4 FILLER_0_41_243 ();
 sg13g2_fill_1 FILLER_0_41_247 ();
 sg13g2_fill_4 FILLER_0_41_252 ();
 sg13g2_fill_4 FILLER_0_41_260 ();
 sg13g2_fill_1 FILLER_0_41_264 ();
 sg13g2_fill_4 FILLER_0_41_269 ();
 sg13g2_fill_1 FILLER_0_41_273 ();
 sg13g2_fill_4 FILLER_0_41_278 ();
 sg13g2_fill_1 FILLER_0_41_282 ();
 sg13g2_fill_2 FILLER_0_41_287 ();
 sg13g2_fill_8 FILLER_0_41_292 ();
 sg13g2_fill_8 FILLER_0_41_300 ();
 sg13g2_fill_4 FILLER_0_41_308 ();
 sg13g2_fill_2 FILLER_0_41_320 ();
 sg13g2_fill_1 FILLER_0_41_322 ();
 sg13g2_fill_2 FILLER_0_42_0 ();
 sg13g2_fill_4 FILLER_0_42_6 ();
 sg13g2_fill_4 FILLER_0_42_14 ();
 sg13g2_fill_1 FILLER_0_42_18 ();
 sg13g2_fill_2 FILLER_0_42_23 ();
 sg13g2_fill_2 FILLER_0_42_33 ();
 sg13g2_fill_2 FILLER_0_42_61 ();
 sg13g2_fill_1 FILLER_0_42_63 ();
 sg13g2_fill_2 FILLER_0_42_90 ();
 sg13g2_fill_4 FILLER_0_42_97 ();
 sg13g2_fill_2 FILLER_0_42_106 ();
 sg13g2_fill_2 FILLER_0_42_134 ();
 sg13g2_fill_1 FILLER_0_42_136 ();
 sg13g2_fill_4 FILLER_0_42_141 ();
 sg13g2_fill_2 FILLER_0_42_150 ();
 sg13g2_fill_1 FILLER_0_42_152 ();
 sg13g2_fill_4 FILLER_0_42_159 ();
 sg13g2_fill_2 FILLER_0_42_189 ();
 sg13g2_fill_1 FILLER_0_42_191 ();
 sg13g2_fill_2 FILLER_0_42_198 ();
 sg13g2_fill_1 FILLER_0_42_200 ();
 sg13g2_fill_2 FILLER_0_42_206 ();
 sg13g2_fill_2 FILLER_0_42_213 ();
 sg13g2_fill_2 FILLER_0_42_221 ();
 sg13g2_fill_1 FILLER_0_42_223 ();
 sg13g2_fill_2 FILLER_0_42_232 ();
 sg13g2_fill_1 FILLER_0_42_234 ();
 sg13g2_fill_4 FILLER_0_42_240 ();
 sg13g2_fill_2 FILLER_0_42_244 ();
 sg13g2_fill_2 FILLER_0_42_251 ();
 sg13g2_fill_2 FILLER_0_42_259 ();
 sg13g2_fill_4 FILLER_0_42_269 ();
 sg13g2_fill_1 FILLER_0_42_273 ();
 sg13g2_fill_2 FILLER_0_42_280 ();
 sg13g2_fill_8 FILLER_0_42_287 ();
 sg13g2_fill_2 FILLER_0_42_321 ();
 sg13g2_fill_1 FILLER_0_43_0 ();
 sg13g2_fill_2 FILLER_0_43_5 ();
 sg13g2_fill_2 FILLER_0_43_11 ();
 sg13g2_fill_2 FILLER_0_43_17 ();
 sg13g2_fill_2 FILLER_0_43_23 ();
 sg13g2_fill_1 FILLER_0_43_25 ();
 sg13g2_fill_2 FILLER_0_43_30 ();
 sg13g2_fill_2 FILLER_0_43_36 ();
 sg13g2_fill_2 FILLER_0_43_42 ();
 sg13g2_fill_1 FILLER_0_43_44 ();
 sg13g2_fill_4 FILLER_0_43_71 ();
 sg13g2_fill_2 FILLER_0_43_75 ();
 sg13g2_fill_2 FILLER_0_43_82 ();
 sg13g2_fill_2 FILLER_0_43_92 ();
 sg13g2_fill_1 FILLER_0_43_94 ();
 sg13g2_fill_2 FILLER_0_43_101 ();
 sg13g2_fill_2 FILLER_0_43_107 ();
 sg13g2_fill_2 FILLER_0_43_117 ();
 sg13g2_fill_1 FILLER_0_43_119 ();
 sg13g2_fill_4 FILLER_0_43_125 ();
 sg13g2_fill_2 FILLER_0_43_134 ();
 sg13g2_fill_1 FILLER_0_43_136 ();
 sg13g2_fill_4 FILLER_0_43_141 ();
 sg13g2_fill_8 FILLER_0_43_150 ();
 sg13g2_fill_4 FILLER_0_43_158 ();
 sg13g2_fill_1 FILLER_0_43_162 ();
 sg13g2_fill_2 FILLER_0_43_170 ();
 sg13g2_fill_4 FILLER_0_43_176 ();
 sg13g2_fill_2 FILLER_0_43_185 ();
 sg13g2_fill_1 FILLER_0_43_187 ();
 sg13g2_fill_4 FILLER_0_43_195 ();
 sg13g2_fill_1 FILLER_0_43_199 ();
 sg13g2_fill_2 FILLER_0_43_204 ();
 sg13g2_fill_2 FILLER_0_43_212 ();
 sg13g2_fill_2 FILLER_0_43_224 ();
 sg13g2_fill_2 FILLER_0_43_234 ();
 sg13g2_fill_2 FILLER_0_43_246 ();
 sg13g2_fill_2 FILLER_0_43_253 ();
 sg13g2_fill_2 FILLER_0_43_259 ();
 sg13g2_fill_8 FILLER_0_43_265 ();
 sg13g2_fill_1 FILLER_0_43_273 ();
 sg13g2_fill_2 FILLER_0_43_279 ();
 sg13g2_fill_2 FILLER_0_43_285 ();
 sg13g2_fill_2 FILLER_0_43_292 ();
 sg13g2_fill_4 FILLER_0_43_298 ();
 sg13g2_fill_2 FILLER_0_43_306 ();
 sg13g2_fill_8 FILLER_0_43_314 ();
 sg13g2_fill_1 FILLER_0_43_322 ();
 sg13g2_fill_2 FILLER_0_44_0 ();
 sg13g2_fill_1 FILLER_0_44_2 ();
 sg13g2_fill_4 FILLER_0_44_29 ();
 sg13g2_fill_2 FILLER_0_44_33 ();
 sg13g2_fill_1 FILLER_0_44_35 ();
 sg13g2_fill_2 FILLER_0_44_44 ();
 sg13g2_fill_1 FILLER_0_44_46 ();
 sg13g2_fill_4 FILLER_0_44_73 ();
 sg13g2_fill_1 FILLER_0_44_77 ();
 sg13g2_fill_2 FILLER_0_44_86 ();
 sg13g2_fill_2 FILLER_0_44_93 ();
 sg13g2_fill_2 FILLER_0_44_99 ();
 sg13g2_fill_1 FILLER_0_44_101 ();
 sg13g2_fill_4 FILLER_0_44_107 ();
 sg13g2_fill_4 FILLER_0_44_119 ();
 sg13g2_fill_2 FILLER_0_44_123 ();
 sg13g2_fill_2 FILLER_0_44_129 ();
 sg13g2_fill_1 FILLER_0_44_131 ();
 sg13g2_fill_2 FILLER_0_44_140 ();
 sg13g2_fill_2 FILLER_0_44_146 ();
 sg13g2_fill_2 FILLER_0_44_153 ();
 sg13g2_fill_2 FILLER_0_44_161 ();
 sg13g2_fill_2 FILLER_0_44_168 ();
 sg13g2_fill_4 FILLER_0_44_175 ();
 sg13g2_fill_2 FILLER_0_44_187 ();
 sg13g2_fill_1 FILLER_0_44_189 ();
 sg13g2_fill_2 FILLER_0_44_194 ();
 sg13g2_fill_2 FILLER_0_44_203 ();
 sg13g2_fill_2 FILLER_0_44_211 ();
 sg13g2_fill_2 FILLER_0_44_218 ();
 sg13g2_fill_4 FILLER_0_44_225 ();
 sg13g2_fill_2 FILLER_0_44_235 ();
 sg13g2_fill_2 FILLER_0_44_242 ();
 sg13g2_fill_2 FILLER_0_44_270 ();
 sg13g2_fill_1 FILLER_0_44_272 ();
 sg13g2_fill_2 FILLER_0_44_279 ();
 sg13g2_fill_4 FILLER_0_44_286 ();
 sg13g2_fill_2 FILLER_0_44_298 ();
 sg13g2_fill_2 FILLER_0_44_308 ();
 sg13g2_fill_8 FILLER_0_44_314 ();
 sg13g2_fill_1 FILLER_0_44_322 ();
 sg13g2_fill_2 FILLER_0_45_0 ();
 sg13g2_fill_1 FILLER_0_45_2 ();
 sg13g2_fill_2 FILLER_0_45_29 ();
 sg13g2_fill_2 FILLER_0_45_36 ();
 sg13g2_fill_4 FILLER_0_45_44 ();
 sg13g2_fill_4 FILLER_0_45_52 ();
 sg13g2_fill_2 FILLER_0_45_56 ();
 sg13g2_fill_1 FILLER_0_45_58 ();
 sg13g2_fill_2 FILLER_0_45_64 ();
 sg13g2_fill_1 FILLER_0_45_66 ();
 sg13g2_fill_4 FILLER_0_45_93 ();
 sg13g2_fill_2 FILLER_0_45_123 ();
 sg13g2_fill_1 FILLER_0_45_125 ();
 sg13g2_fill_2 FILLER_0_45_131 ();
 sg13g2_fill_1 FILLER_0_45_133 ();
 sg13g2_fill_4 FILLER_0_45_140 ();
 sg13g2_fill_4 FILLER_0_45_149 ();
 sg13g2_fill_4 FILLER_0_45_158 ();
 sg13g2_fill_1 FILLER_0_45_162 ();
 sg13g2_fill_4 FILLER_0_45_167 ();
 sg13g2_fill_4 FILLER_0_45_179 ();
 sg13g2_fill_1 FILLER_0_45_183 ();
 sg13g2_fill_2 FILLER_0_45_191 ();
 sg13g2_fill_1 FILLER_0_45_193 ();
 sg13g2_fill_2 FILLER_0_45_199 ();
 sg13g2_fill_2 FILLER_0_45_211 ();
 sg13g2_fill_1 FILLER_0_45_213 ();
 sg13g2_fill_4 FILLER_0_45_222 ();
 sg13g2_fill_2 FILLER_0_45_226 ();
 sg13g2_fill_2 FILLER_0_45_233 ();
 sg13g2_fill_8 FILLER_0_45_261 ();
 sg13g2_fill_1 FILLER_0_45_269 ();
 sg13g2_fill_2 FILLER_0_45_273 ();
 sg13g2_fill_4 FILLER_0_45_280 ();
 sg13g2_fill_4 FILLER_0_45_288 ();
 sg13g2_fill_1 FILLER_0_45_292 ();
 sg13g2_fill_2 FILLER_0_45_297 ();
 sg13g2_fill_4 FILLER_0_45_304 ();
 sg13g2_fill_2 FILLER_0_45_308 ();
 sg13g2_fill_1 FILLER_0_45_310 ();
 sg13g2_fill_4 FILLER_0_45_319 ();
 sg13g2_fill_2 FILLER_0_46_0 ();
 sg13g2_fill_1 FILLER_0_46_2 ();
 sg13g2_fill_2 FILLER_0_46_7 ();
 sg13g2_fill_2 FILLER_0_46_14 ();
 sg13g2_fill_2 FILLER_0_46_20 ();
 sg13g2_fill_2 FILLER_0_46_26 ();
 sg13g2_fill_1 FILLER_0_46_28 ();
 sg13g2_fill_2 FILLER_0_46_37 ();
 sg13g2_fill_1 FILLER_0_46_39 ();
 sg13g2_fill_4 FILLER_0_46_45 ();
 sg13g2_fill_1 FILLER_0_46_49 ();
 sg13g2_fill_2 FILLER_0_46_54 ();
 sg13g2_fill_4 FILLER_0_46_61 ();
 sg13g2_fill_2 FILLER_0_46_65 ();
 sg13g2_fill_1 FILLER_0_46_67 ();
 sg13g2_fill_2 FILLER_0_46_72 ();
 sg13g2_fill_2 FILLER_0_46_78 ();
 sg13g2_fill_4 FILLER_0_46_85 ();
 sg13g2_fill_4 FILLER_0_46_97 ();
 sg13g2_fill_1 FILLER_0_46_101 ();
 sg13g2_fill_4 FILLER_0_46_107 ();
 sg13g2_fill_2 FILLER_0_46_115 ();
 sg13g2_fill_1 FILLER_0_46_117 ();
 sg13g2_fill_4 FILLER_0_46_125 ();
 sg13g2_fill_2 FILLER_0_46_134 ();
 sg13g2_fill_1 FILLER_0_46_136 ();
 sg13g2_fill_2 FILLER_0_46_149 ();
 sg13g2_fill_8 FILLER_0_46_159 ();
 sg13g2_fill_8 FILLER_0_46_167 ();
 sg13g2_fill_8 FILLER_0_46_175 ();
 sg13g2_fill_2 FILLER_0_46_187 ();
 sg13g2_fill_2 FILLER_0_46_194 ();
 sg13g2_fill_4 FILLER_0_46_201 ();
 sg13g2_fill_2 FILLER_0_46_205 ();
 sg13g2_fill_4 FILLER_0_46_212 ();
 sg13g2_fill_2 FILLER_0_46_221 ();
 sg13g2_fill_2 FILLER_0_46_227 ();
 sg13g2_fill_2 FILLER_0_46_237 ();
 sg13g2_fill_2 FILLER_0_46_265 ();
 sg13g2_fill_2 FILLER_0_46_270 ();
 sg13g2_fill_2 FILLER_0_46_277 ();
 sg13g2_fill_1 FILLER_0_46_279 ();
 sg13g2_fill_2 FILLER_0_46_285 ();
 sg13g2_fill_2 FILLER_0_46_293 ();
 sg13g2_fill_2 FILLER_0_46_321 ();
 sg13g2_fill_2 FILLER_0_47_0 ();
 sg13g2_fill_2 FILLER_0_47_7 ();
 sg13g2_fill_2 FILLER_0_47_14 ();
 sg13g2_fill_2 FILLER_0_47_21 ();
 sg13g2_fill_2 FILLER_0_47_26 ();
 sg13g2_fill_2 FILLER_0_47_31 ();
 sg13g2_fill_2 FILLER_0_47_37 ();
 sg13g2_fill_2 FILLER_0_47_65 ();
 sg13g2_fill_2 FILLER_0_47_71 ();
 sg13g2_fill_2 FILLER_0_47_99 ();
 sg13g2_fill_2 FILLER_0_47_104 ();
 sg13g2_fill_2 FILLER_0_47_132 ();
 sg13g2_fill_2 FILLER_0_47_143 ();
 sg13g2_fill_2 FILLER_0_47_151 ();
 sg13g2_fill_2 FILLER_0_47_157 ();
 sg13g2_fill_8 FILLER_0_47_164 ();
 sg13g2_fill_2 FILLER_0_47_172 ();
 sg13g2_fill_2 FILLER_0_47_179 ();
 sg13g2_fill_1 FILLER_0_47_181 ();
 sg13g2_fill_4 FILLER_0_47_187 ();
 sg13g2_fill_2 FILLER_0_47_195 ();
 sg13g2_fill_4 FILLER_0_47_202 ();
 sg13g2_fill_2 FILLER_0_47_212 ();
 sg13g2_fill_4 FILLER_0_47_219 ();
 sg13g2_fill_2 FILLER_0_47_223 ();
 sg13g2_fill_1 FILLER_0_47_225 ();
 sg13g2_fill_2 FILLER_0_47_232 ();
 sg13g2_fill_2 FILLER_0_47_239 ();
 sg13g2_fill_4 FILLER_0_47_246 ();
 sg13g2_fill_1 FILLER_0_47_250 ();
 sg13g2_fill_4 FILLER_0_47_256 ();
 sg13g2_fill_4 FILLER_0_47_268 ();
 sg13g2_fill_2 FILLER_0_47_272 ();
 sg13g2_fill_1 FILLER_0_47_274 ();
 sg13g2_fill_2 FILLER_0_47_281 ();
 sg13g2_fill_4 FILLER_0_47_288 ();
 sg13g2_fill_4 FILLER_0_47_296 ();
 sg13g2_fill_4 FILLER_0_47_308 ();
 sg13g2_fill_2 FILLER_0_47_320 ();
 sg13g2_fill_1 FILLER_0_47_322 ();
 sg13g2_fill_4 FILLER_0_48_0 ();
 sg13g2_fill_2 FILLER_0_48_4 ();
 sg13g2_fill_2 FILLER_0_48_11 ();
 sg13g2_fill_2 FILLER_0_48_18 ();
 sg13g2_fill_2 FILLER_0_48_24 ();
 sg13g2_fill_4 FILLER_0_48_38 ();
 sg13g2_fill_1 FILLER_0_48_42 ();
 sg13g2_fill_2 FILLER_0_48_47 ();
 sg13g2_fill_4 FILLER_0_48_53 ();
 sg13g2_fill_4 FILLER_0_48_62 ();
 sg13g2_fill_1 FILLER_0_48_66 ();
 sg13g2_fill_4 FILLER_0_48_71 ();
 sg13g2_fill_1 FILLER_0_48_75 ();
 sg13g2_fill_4 FILLER_0_48_84 ();
 sg13g2_fill_1 FILLER_0_48_88 ();
 sg13g2_fill_2 FILLER_0_48_94 ();
 sg13g2_fill_2 FILLER_0_48_101 ();
 sg13g2_fill_4 FILLER_0_48_129 ();
 sg13g2_fill_2 FILLER_0_48_136 ();
 sg13g2_fill_4 FILLER_0_48_142 ();
 sg13g2_fill_4 FILLER_0_48_154 ();
 sg13g2_fill_1 FILLER_0_48_158 ();
 sg13g2_fill_8 FILLER_0_48_163 ();
 sg13g2_fill_2 FILLER_0_48_171 ();
 sg13g2_fill_4 FILLER_0_48_178 ();
 sg13g2_fill_2 FILLER_0_48_182 ();
 sg13g2_fill_4 FILLER_0_48_189 ();
 sg13g2_fill_4 FILLER_0_48_199 ();
 sg13g2_fill_1 FILLER_0_48_203 ();
 sg13g2_fill_2 FILLER_0_48_212 ();
 sg13g2_fill_4 FILLER_0_48_220 ();
 sg13g2_fill_2 FILLER_0_48_228 ();
 sg13g2_fill_2 FILLER_0_48_256 ();
 sg13g2_fill_8 FILLER_0_48_284 ();
 sg13g2_fill_4 FILLER_0_48_292 ();
 sg13g2_fill_2 FILLER_0_48_296 ();
 sg13g2_fill_2 FILLER_0_48_302 ();
 sg13g2_fill_2 FILLER_0_48_308 ();
 sg13g2_fill_4 FILLER_0_48_318 ();
 sg13g2_fill_1 FILLER_0_48_322 ();
 sg13g2_fill_2 FILLER_0_49_0 ();
 sg13g2_fill_2 FILLER_0_49_28 ();
 sg13g2_fill_1 FILLER_0_49_30 ();
 sg13g2_fill_2 FILLER_0_49_36 ();
 sg13g2_fill_2 FILLER_0_49_44 ();
 sg13g2_fill_2 FILLER_0_49_52 ();
 sg13g2_fill_2 FILLER_0_49_59 ();
 sg13g2_fill_1 FILLER_0_49_61 ();
 sg13g2_fill_2 FILLER_0_49_67 ();
 sg13g2_fill_2 FILLER_0_49_72 ();
 sg13g2_fill_1 FILLER_0_49_74 ();
 sg13g2_fill_4 FILLER_0_49_79 ();
 sg13g2_fill_2 FILLER_0_49_83 ();
 sg13g2_fill_2 FILLER_0_49_90 ();
 sg13g2_fill_4 FILLER_0_49_95 ();
 sg13g2_fill_2 FILLER_0_49_99 ();
 sg13g2_fill_2 FILLER_0_49_106 ();
 sg13g2_fill_4 FILLER_0_49_112 ();
 sg13g2_fill_2 FILLER_0_49_116 ();
 sg13g2_fill_2 FILLER_0_49_126 ();
 sg13g2_fill_1 FILLER_0_49_128 ();
 sg13g2_fill_2 FILLER_0_49_133 ();
 sg13g2_fill_8 FILLER_0_49_140 ();
 sg13g2_fill_8 FILLER_0_49_148 ();
 sg13g2_fill_1 FILLER_0_49_156 ();
 sg13g2_fill_8 FILLER_0_49_160 ();
 sg13g2_fill_2 FILLER_0_49_168 ();
 sg13g2_fill_1 FILLER_0_49_170 ();
 sg13g2_fill_2 FILLER_0_49_176 ();
 sg13g2_fill_4 FILLER_0_49_182 ();
 sg13g2_fill_2 FILLER_0_49_186 ();
 sg13g2_fill_1 FILLER_0_49_188 ();
 sg13g2_fill_2 FILLER_0_49_193 ();
 sg13g2_fill_1 FILLER_0_49_195 ();
 sg13g2_fill_2 FILLER_0_49_200 ();
 sg13g2_fill_2 FILLER_0_49_208 ();
 sg13g2_fill_2 FILLER_0_49_215 ();
 sg13g2_fill_8 FILLER_0_49_222 ();
 sg13g2_fill_8 FILLER_0_49_230 ();
 sg13g2_fill_4 FILLER_0_49_238 ();
 sg13g2_fill_1 FILLER_0_49_242 ();
 sg13g2_fill_2 FILLER_0_49_247 ();
 sg13g2_fill_2 FILLER_0_49_253 ();
 sg13g2_fill_2 FILLER_0_49_259 ();
 sg13g2_fill_2 FILLER_0_49_265 ();
 sg13g2_fill_4 FILLER_0_49_271 ();
 sg13g2_fill_2 FILLER_0_49_275 ();
 sg13g2_fill_2 FILLER_0_49_284 ();
 sg13g2_fill_2 FILLER_0_49_290 ();
 sg13g2_fill_2 FILLER_0_49_297 ();
 sg13g2_fill_4 FILLER_0_49_304 ();
 sg13g2_fill_2 FILLER_0_49_308 ();
 sg13g2_fill_1 FILLER_0_49_310 ();
 sg13g2_fill_2 FILLER_0_49_316 ();
 sg13g2_fill_1 FILLER_0_49_322 ();
 sg13g2_fill_2 FILLER_0_50_0 ();
 sg13g2_fill_2 FILLER_0_50_6 ();
 sg13g2_fill_1 FILLER_0_50_8 ();
 sg13g2_fill_2 FILLER_0_50_13 ();
 sg13g2_fill_1 FILLER_0_50_15 ();
 sg13g2_fill_4 FILLER_0_50_20 ();
 sg13g2_fill_2 FILLER_0_50_27 ();
 sg13g2_fill_1 FILLER_0_50_29 ();
 sg13g2_fill_2 FILLER_0_50_35 ();
 sg13g2_fill_2 FILLER_0_50_41 ();
 sg13g2_fill_1 FILLER_0_50_43 ();
 sg13g2_fill_2 FILLER_0_50_50 ();
 sg13g2_fill_2 FILLER_0_50_56 ();
 sg13g2_fill_2 FILLER_0_50_63 ();
 sg13g2_fill_2 FILLER_0_50_70 ();
 sg13g2_fill_2 FILLER_0_50_80 ();
 sg13g2_fill_8 FILLER_0_50_87 ();
 sg13g2_fill_2 FILLER_0_50_95 ();
 sg13g2_fill_1 FILLER_0_50_97 ();
 sg13g2_fill_4 FILLER_0_50_106 ();
 sg13g2_fill_2 FILLER_0_50_110 ();
 sg13g2_fill_1 FILLER_0_50_112 ();
 sg13g2_fill_4 FILLER_0_50_117 ();
 sg13g2_fill_2 FILLER_0_50_121 ();
 sg13g2_fill_1 FILLER_0_50_123 ();
 sg13g2_fill_2 FILLER_0_50_132 ();
 sg13g2_fill_1 FILLER_0_50_134 ();
 sg13g2_fill_2 FILLER_0_50_143 ();
 sg13g2_fill_1 FILLER_0_50_145 ();
 sg13g2_fill_4 FILLER_0_50_150 ();
 sg13g2_fill_2 FILLER_0_50_158 ();
 sg13g2_fill_1 FILLER_0_50_160 ();
 sg13g2_fill_4 FILLER_0_50_165 ();
 sg13g2_fill_2 FILLER_0_50_176 ();
 sg13g2_fill_1 FILLER_0_50_178 ();
 sg13g2_fill_2 FILLER_0_50_185 ();
 sg13g2_fill_8 FILLER_0_50_192 ();
 sg13g2_fill_1 FILLER_0_50_200 ();
 sg13g2_fill_2 FILLER_0_50_206 ();
 sg13g2_fill_2 FILLER_0_50_216 ();
 sg13g2_fill_2 FILLER_0_50_223 ();
 sg13g2_fill_1 FILLER_0_50_225 ();
 sg13g2_fill_2 FILLER_0_50_232 ();
 sg13g2_fill_1 FILLER_0_50_234 ();
 sg13g2_fill_2 FILLER_0_50_239 ();
 sg13g2_fill_1 FILLER_0_50_241 ();
 sg13g2_fill_2 FILLER_0_50_247 ();
 sg13g2_fill_1 FILLER_0_50_249 ();
 sg13g2_fill_2 FILLER_0_50_253 ();
 sg13g2_fill_1 FILLER_0_50_255 ();
 sg13g2_fill_2 FILLER_0_50_262 ();
 sg13g2_fill_1 FILLER_0_50_264 ();
 sg13g2_fill_2 FILLER_0_50_270 ();
 sg13g2_fill_4 FILLER_0_50_276 ();
 sg13g2_fill_2 FILLER_0_50_288 ();
 sg13g2_fill_2 FILLER_0_50_295 ();
 sg13g2_fill_2 FILLER_0_50_305 ();
 sg13g2_fill_1 FILLER_0_50_307 ();
 sg13g2_fill_2 FILLER_0_50_314 ();
 sg13g2_fill_2 FILLER_0_50_320 ();
 sg13g2_fill_1 FILLER_0_50_322 ();
 sg13g2_fill_2 FILLER_0_51_0 ();
 sg13g2_fill_2 FILLER_0_51_28 ();
 sg13g2_fill_2 FILLER_0_51_38 ();
 sg13g2_fill_2 FILLER_0_51_44 ();
 sg13g2_fill_2 FILLER_0_51_49 ();
 sg13g2_fill_2 FILLER_0_51_55 ();
 sg13g2_fill_2 FILLER_0_51_61 ();
 sg13g2_fill_2 FILLER_0_51_68 ();
 sg13g2_fill_2 FILLER_0_51_74 ();
 sg13g2_fill_2 FILLER_0_51_81 ();
 sg13g2_fill_2 FILLER_0_51_109 ();
 sg13g2_fill_2 FILLER_0_51_115 ();
 sg13g2_fill_1 FILLER_0_51_117 ();
 sg13g2_fill_2 FILLER_0_51_123 ();
 sg13g2_fill_1 FILLER_0_51_125 ();
 sg13g2_fill_2 FILLER_0_51_152 ();
 sg13g2_fill_2 FILLER_0_51_158 ();
 sg13g2_fill_1 FILLER_0_51_160 ();
 sg13g2_fill_2 FILLER_0_51_166 ();
 sg13g2_fill_2 FILLER_0_51_174 ();
 sg13g2_fill_4 FILLER_0_51_182 ();
 sg13g2_fill_2 FILLER_0_51_189 ();
 sg13g2_fill_8 FILLER_0_51_198 ();
 sg13g2_fill_4 FILLER_0_51_206 ();
 sg13g2_fill_2 FILLER_0_51_210 ();
 sg13g2_fill_2 FILLER_0_51_216 ();
 sg13g2_fill_1 FILLER_0_51_218 ();
 sg13g2_fill_4 FILLER_0_51_224 ();
 sg13g2_fill_4 FILLER_0_51_254 ();
 sg13g2_fill_4 FILLER_0_51_262 ();
 sg13g2_fill_2 FILLER_0_51_274 ();
 sg13g2_fill_2 FILLER_0_51_280 ();
 sg13g2_fill_2 FILLER_0_51_287 ();
 sg13g2_fill_2 FILLER_0_51_295 ();
 sg13g2_fill_4 FILLER_0_51_305 ();
 sg13g2_fill_2 FILLER_0_51_315 ();
 sg13g2_fill_2 FILLER_0_51_321 ();
 sg13g2_fill_4 FILLER_0_52_0 ();
 sg13g2_fill_2 FILLER_0_52_30 ();
 sg13g2_fill_2 FILLER_0_52_36 ();
 sg13g2_fill_1 FILLER_0_52_38 ();
 sg13g2_fill_2 FILLER_0_52_43 ();
 sg13g2_fill_1 FILLER_0_52_45 ();
 sg13g2_fill_4 FILLER_0_52_51 ();
 sg13g2_fill_2 FILLER_0_52_59 ();
 sg13g2_fill_2 FILLER_0_52_66 ();
 sg13g2_fill_2 FILLER_0_52_76 ();
 sg13g2_fill_4 FILLER_0_52_82 ();
 sg13g2_fill_1 FILLER_0_52_86 ();
 sg13g2_fill_2 FILLER_0_52_95 ();
 sg13g2_fill_4 FILLER_0_52_123 ();
 sg13g2_fill_1 FILLER_0_52_127 ();
 sg13g2_fill_2 FILLER_0_52_154 ();
 sg13g2_fill_1 FILLER_0_52_156 ();
 sg13g2_fill_2 FILLER_0_52_161 ();
 sg13g2_fill_2 FILLER_0_52_168 ();
 sg13g2_fill_2 FILLER_0_52_175 ();
 sg13g2_fill_2 FILLER_0_52_183 ();
 sg13g2_fill_4 FILLER_0_52_190 ();
 sg13g2_fill_8 FILLER_0_52_199 ();
 sg13g2_fill_8 FILLER_0_52_207 ();
 sg13g2_fill_1 FILLER_0_52_215 ();
 sg13g2_fill_4 FILLER_0_52_220 ();
 sg13g2_fill_2 FILLER_0_52_229 ();
 sg13g2_fill_1 FILLER_0_52_231 ();
 sg13g2_fill_2 FILLER_0_52_258 ();
 sg13g2_fill_4 FILLER_0_52_286 ();
 sg13g2_fill_2 FILLER_0_52_290 ();
 sg13g2_fill_2 FILLER_0_52_297 ();
 sg13g2_fill_2 FILLER_0_52_302 ();
 sg13g2_fill_2 FILLER_0_52_312 ();
 sg13g2_fill_4 FILLER_0_52_318 ();
 sg13g2_fill_1 FILLER_0_52_322 ();
 sg13g2_fill_2 FILLER_0_53_0 ();
 sg13g2_fill_4 FILLER_0_53_6 ();
 sg13g2_fill_2 FILLER_0_53_14 ();
 sg13g2_fill_1 FILLER_0_53_16 ();
 sg13g2_fill_4 FILLER_0_53_25 ();
 sg13g2_fill_2 FILLER_0_53_34 ();
 sg13g2_fill_1 FILLER_0_53_36 ();
 sg13g2_fill_4 FILLER_0_53_42 ();
 sg13g2_fill_2 FILLER_0_53_50 ();
 sg13g2_fill_4 FILLER_0_53_55 ();
 sg13g2_fill_2 FILLER_0_53_59 ();
 sg13g2_fill_1 FILLER_0_53_61 ();
 sg13g2_fill_2 FILLER_0_53_66 ();
 sg13g2_fill_1 FILLER_0_53_68 ();
 sg13g2_fill_2 FILLER_0_53_76 ();
 sg13g2_fill_1 FILLER_0_53_78 ();
 sg13g2_fill_4 FILLER_0_53_83 ();
 sg13g2_fill_1 FILLER_0_53_87 ();
 sg13g2_fill_2 FILLER_0_53_92 ();
 sg13g2_fill_2 FILLER_0_53_98 ();
 sg13g2_fill_4 FILLER_0_53_104 ();
 sg13g2_fill_2 FILLER_0_53_116 ();
 sg13g2_fill_1 FILLER_0_53_118 ();
 sg13g2_fill_2 FILLER_0_53_123 ();
 sg13g2_fill_2 FILLER_0_53_130 ();
 sg13g2_fill_1 FILLER_0_53_132 ();
 sg13g2_fill_2 FILLER_0_53_136 ();
 sg13g2_fill_2 FILLER_0_53_142 ();
 sg13g2_fill_2 FILLER_0_53_152 ();
 sg13g2_fill_8 FILLER_0_53_158 ();
 sg13g2_fill_2 FILLER_0_53_172 ();
 sg13g2_fill_2 FILLER_0_53_179 ();
 sg13g2_fill_2 FILLER_0_53_186 ();
 sg13g2_fill_2 FILLER_0_53_192 ();
 sg13g2_fill_4 FILLER_0_53_199 ();
 sg13g2_fill_2 FILLER_0_53_207 ();
 sg13g2_fill_2 FILLER_0_53_214 ();
 sg13g2_fill_2 FILLER_0_53_221 ();
 sg13g2_fill_2 FILLER_0_53_227 ();
 sg13g2_fill_2 FILLER_0_53_233 ();
 sg13g2_fill_2 FILLER_0_53_261 ();
 sg13g2_fill_2 FILLER_0_53_271 ();
 sg13g2_fill_2 FILLER_0_53_277 ();
 sg13g2_fill_2 FILLER_0_53_286 ();
 sg13g2_fill_2 FILLER_0_53_296 ();
 sg13g2_fill_2 FILLER_0_53_302 ();
 sg13g2_fill_2 FILLER_0_53_312 ();
 sg13g2_fill_1 FILLER_0_53_322 ();
 sg13g2_fill_4 FILLER_0_54_0 ();
 sg13g2_fill_2 FILLER_0_54_4 ();
 sg13g2_fill_1 FILLER_0_54_6 ();
 sg13g2_fill_2 FILLER_0_54_11 ();
 sg13g2_fill_2 FILLER_0_54_17 ();
 sg13g2_fill_4 FILLER_0_54_23 ();
 sg13g2_fill_2 FILLER_0_54_32 ();
 sg13g2_fill_2 FILLER_0_54_39 ();
 sg13g2_fill_2 FILLER_0_54_46 ();
 sg13g2_fill_2 FILLER_0_54_52 ();
 sg13g2_fill_2 FILLER_0_54_59 ();
 sg13g2_fill_2 FILLER_0_54_66 ();
 sg13g2_fill_4 FILLER_0_54_73 ();
 sg13g2_fill_2 FILLER_0_54_85 ();
 sg13g2_fill_2 FILLER_0_54_113 ();
 sg13g2_fill_2 FILLER_0_54_141 ();
 sg13g2_fill_2 FILLER_0_54_147 ();
 sg13g2_fill_1 FILLER_0_54_149 ();
 sg13g2_fill_2 FILLER_0_54_176 ();
 sg13g2_fill_2 FILLER_0_54_182 ();
 sg13g2_fill_1 FILLER_0_54_184 ();
 sg13g2_fill_4 FILLER_0_54_191 ();
 sg13g2_fill_2 FILLER_0_54_221 ();
 sg13g2_fill_1 FILLER_0_54_223 ();
 sg13g2_fill_4 FILLER_0_54_228 ();
 sg13g2_fill_2 FILLER_0_54_236 ();
 sg13g2_fill_2 FILLER_0_54_242 ();
 sg13g2_fill_4 FILLER_0_54_248 ();
 sg13g2_fill_2 FILLER_0_54_257 ();
 sg13g2_fill_2 FILLER_0_54_265 ();
 sg13g2_fill_1 FILLER_0_54_267 ();
 sg13g2_fill_2 FILLER_0_54_272 ();
 sg13g2_fill_4 FILLER_0_54_282 ();
 sg13g2_fill_1 FILLER_0_54_286 ();
 sg13g2_fill_2 FILLER_0_54_291 ();
 sg13g2_fill_2 FILLER_0_54_301 ();
 sg13g2_fill_4 FILLER_0_54_307 ();
 sg13g2_fill_8 FILLER_0_54_315 ();
 sg13g2_fill_2 FILLER_0_55_0 ();
 sg13g2_fill_1 FILLER_0_55_2 ();
 sg13g2_fill_2 FILLER_0_55_7 ();
 sg13g2_fill_2 FILLER_0_55_12 ();
 sg13g2_fill_1 FILLER_0_55_14 ();
 sg13g2_fill_2 FILLER_0_55_19 ();
 sg13g2_fill_2 FILLER_0_55_47 ();
 sg13g2_fill_1 FILLER_0_55_49 ();
 sg13g2_fill_4 FILLER_0_55_55 ();
 sg13g2_fill_2 FILLER_0_55_59 ();
 sg13g2_fill_2 FILLER_0_55_66 ();
 sg13g2_fill_8 FILLER_0_55_76 ();
 sg13g2_fill_4 FILLER_0_55_84 ();
 sg13g2_fill_1 FILLER_0_55_88 ();
 sg13g2_fill_2 FILLER_0_55_97 ();
 sg13g2_fill_1 FILLER_0_55_99 ();
 sg13g2_fill_2 FILLER_0_55_104 ();
 sg13g2_fill_2 FILLER_0_55_132 ();
 sg13g2_fill_1 FILLER_0_55_134 ();
 sg13g2_fill_2 FILLER_0_55_161 ();
 sg13g2_fill_1 FILLER_0_55_163 ();
 sg13g2_fill_4 FILLER_0_55_168 ();
 sg13g2_fill_4 FILLER_0_55_177 ();
 sg13g2_fill_2 FILLER_0_55_185 ();
 sg13g2_fill_1 FILLER_0_55_187 ();
 sg13g2_fill_2 FILLER_0_55_214 ();
 sg13g2_fill_1 FILLER_0_55_216 ();
 sg13g2_fill_8 FILLER_0_55_243 ();
 sg13g2_fill_2 FILLER_0_55_251 ();
 sg13g2_fill_1 FILLER_0_55_253 ();
 sg13g2_fill_2 FILLER_0_55_261 ();
 sg13g2_fill_2 FILLER_0_55_271 ();
 sg13g2_fill_4 FILLER_0_55_278 ();
 sg13g2_fill_2 FILLER_0_55_282 ();
 sg13g2_fill_1 FILLER_0_55_284 ();
 sg13g2_fill_2 FILLER_0_55_293 ();
 sg13g2_fill_2 FILLER_0_55_321 ();
 sg13g2_fill_4 FILLER_0_56_0 ();
 sg13g2_fill_1 FILLER_0_56_4 ();
 sg13g2_fill_2 FILLER_0_56_31 ();
 sg13g2_fill_2 FILLER_0_56_59 ();
 sg13g2_fill_1 FILLER_0_56_61 ();
 sg13g2_fill_2 FILLER_0_56_66 ();
 sg13g2_fill_2 FILLER_0_56_76 ();
 sg13g2_fill_2 FILLER_0_56_82 ();
 sg13g2_fill_4 FILLER_0_56_110 ();
 sg13g2_fill_2 FILLER_0_56_118 ();
 sg13g2_fill_2 FILLER_0_56_124 ();
 sg13g2_fill_2 FILLER_0_56_152 ();
 sg13g2_fill_1 FILLER_0_56_154 ();
 sg13g2_fill_4 FILLER_0_56_181 ();
 sg13g2_fill_2 FILLER_0_56_185 ();
 sg13g2_fill_2 FILLER_0_56_213 ();
 sg13g2_fill_2 FILLER_0_56_241 ();
 sg13g2_fill_1 FILLER_0_56_243 ();
 sg13g2_fill_2 FILLER_0_56_252 ();
 sg13g2_fill_2 FILLER_0_56_259 ();
 sg13g2_fill_4 FILLER_0_56_265 ();
 sg13g2_fill_2 FILLER_0_56_277 ();
 sg13g2_fill_1 FILLER_0_56_279 ();
 sg13g2_fill_4 FILLER_0_56_306 ();
 sg13g2_fill_1 FILLER_0_56_310 ();
 sg13g2_fill_4 FILLER_0_56_319 ();
 sg13g2_fill_4 FILLER_0_57_0 ();
 sg13g2_fill_2 FILLER_0_57_8 ();
 sg13g2_fill_2 FILLER_0_57_14 ();
 sg13g2_fill_2 FILLER_0_57_20 ();
 sg13g2_fill_2 FILLER_0_57_26 ();
 sg13g2_fill_2 FILLER_0_57_32 ();
 sg13g2_fill_2 FILLER_0_57_38 ();
 sg13g2_fill_2 FILLER_0_57_44 ();
 sg13g2_fill_2 FILLER_0_57_50 ();
 sg13g2_fill_2 FILLER_0_57_56 ();
 sg13g2_fill_2 FILLER_0_57_62 ();
 sg13g2_fill_2 FILLER_0_57_68 ();
 sg13g2_fill_2 FILLER_0_57_96 ();
 sg13g2_fill_2 FILLER_0_57_102 ();
 sg13g2_fill_2 FILLER_0_57_108 ();
 sg13g2_fill_1 FILLER_0_57_110 ();
 sg13g2_fill_2 FILLER_0_57_115 ();
 sg13g2_fill_2 FILLER_0_57_121 ();
 sg13g2_fill_2 FILLER_0_57_127 ();
 sg13g2_fill_2 FILLER_0_57_133 ();
 sg13g2_fill_2 FILLER_0_57_139 ();
 sg13g2_fill_4 FILLER_0_57_145 ();
 sg13g2_fill_2 FILLER_0_57_153 ();
 sg13g2_fill_2 FILLER_0_57_159 ();
 sg13g2_fill_2 FILLER_0_57_165 ();
 sg13g2_fill_2 FILLER_0_57_171 ();
 sg13g2_fill_2 FILLER_0_57_177 ();
 sg13g2_fill_2 FILLER_0_57_184 ();
 sg13g2_fill_2 FILLER_0_57_190 ();
 sg13g2_fill_2 FILLER_0_57_197 ();
 sg13g2_fill_2 FILLER_0_57_203 ();
 sg13g2_fill_2 FILLER_0_57_209 ();
 sg13g2_fill_2 FILLER_0_57_215 ();
 sg13g2_fill_4 FILLER_0_57_221 ();
 sg13g2_fill_2 FILLER_0_57_229 ();
 sg13g2_fill_1 FILLER_0_57_231 ();
 sg13g2_fill_2 FILLER_0_57_239 ();
 sg13g2_fill_1 FILLER_0_57_241 ();
 sg13g2_fill_2 FILLER_0_57_252 ();
 sg13g2_fill_2 FILLER_0_57_260 ();
 sg13g2_fill_2 FILLER_0_57_266 ();
 sg13g2_fill_2 FILLER_0_57_273 ();
 sg13g2_fill_2 FILLER_0_57_280 ();
 sg13g2_fill_2 FILLER_0_57_286 ();
 sg13g2_fill_2 FILLER_0_57_292 ();
 sg13g2_fill_1 FILLER_0_57_294 ();
 sg13g2_fill_2 FILLER_0_57_299 ();
 sg13g2_fill_2 FILLER_0_57_305 ();
 sg13g2_fill_2 FILLER_0_57_311 ();
 sg13g2_fill_4 FILLER_0_57_317 ();
 sg13g2_fill_2 FILLER_0_57_321 ();
 assign uio_oe[0] = net90;
 assign uio_oe[7] = net87;
endmodule
